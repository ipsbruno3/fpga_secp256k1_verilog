precomp_x[0] = 256'h79BE667EF9DCBBAC55A06295CE870B07029BFCDB2DCE28D959F2815B16F81798;
precomp_x[1] = 256'hF9308A019258C31049344F85F89D5229B531C845836F99B08601F113BCE036F9;
precomp_x[2] = 256'h2F8BDE4D1A07209355B4A7250A5C5128E88B84BDDC619AB7CBA8D569B240EFE4;
precomp_x[3] = 256'h5CBDF0646E5DB4EAA398F365F2EA7A0E3D419B7E0330E39CE92BDDEDCAC4F9BC;
precomp_x[4] = 256'hACD484E2F0C7F65309AD178A9F559ABDE09796974C57E714C35F110DFC27CCBE;
precomp_x[5] = 256'h774AE7F858A9411E5EF4246B70C65AAC5649980BE5C17891BBEC17895DA008CB;
precomp_x[6] = 256'hF28773C2D975288BC7D1D205C3748651B075FBC6610E58CDDEEDDF8F19405AA8;
precomp_x[7] = 256'hD7924D4F7D43EA965A465AE3095FF41131E5946F3C85F79E44ADBCF8E27E080E;
precomp_x[8] = 256'hDEFDEA4CDB677750A420FEE807EACF21EB9898AE79B9768766E4FAA04A2D4A34;
precomp_x[9] = 256'h2B4EA0A797A443D293EF5CFF444F4979F06ACFEBD7E86D277475656138385B6C;
precomp_x[10] = 256'h352BBF4A4CDD12564F93FA332CE333301D9AD40271F8107181340AEF25BE59D5;
precomp_x[11] = 256'h2FA2104D6B38D11B0230010559879124E42AB8DFEFF5FF29DC9CDADD4ECACC3F;
precomp_x[12] = 256'h9248279B09B4D68DAB21A9B066EDDA83263C3D84E09572E269CA0CD7F5453714;
precomp_x[13] = 256'hDAED4F2BE3A8BF278E70132FB0BEB7522F570E144BF615C07E996D443DEE8729;
precomp_x[14] = 256'hC44D12C7065D812E8ACF28D7CBB19F9011ECD9E9FDF281B0E6A3B5E87D22E7DB;
precomp_x[15] = 256'h6A245BF6DC698504C89A20CFDED60853152B695336C28063B61C65CBD269E6B4;
precomp_x[16] = 256'h1697FFA6FD9DE627C077E3D2FE541084CE13300B0BEC1146F95AE57F0D0BD6A5;
precomp_x[17] = 256'h605BDB019981718B986D0F07E834CB0D9DEB8360FFB7F61DF982345EF27A7479;
precomp_x[18] = 256'h62D14DAB4150BF497402FDC45A215E10DCB01C354959B10CFE31C7E9D87FF33D;
precomp_x[19] = 256'h80C60AD0040F27DADE5B4B06C408E56B2C50E9F56B9B8B425E555C2F86308B6F;
precomp_x[20] = 256'h7A9375AD6167AD54AA74C6348CC54D344CC5DC9487D847049D5EABB0FA03C8FB;
precomp_x[21] = 256'hD528ECD9B696B54C907A9ED045447A79BB408EC39B68DF504BB51F459BC3FFC9;
precomp_x[22] = 256'h049370A4B5F43412EA25F514E8ECDAD05266115E4A7ECB1387231808F8B45963;
precomp_x[23] = 256'h77F230936EE88CBBD73DF930D64702EF881D811E0E1498E2F1C13EB1FC345D74;
precomp_x[24] = 256'hF2DAC991CC4CE4B9EA44887E5C7C0BCE58C80074AB9D4DBAEB28531B7739F530;
precomp_x[25] = 256'h463B3D9F662621FB1B4BE8FBBE2520125A216CDFC9DAE3DEBCBA4850C690D45B;
precomp_x[26] = 256'hF16F804244E46E2A09232D4AFF3B59976B98FAC14328A2D1A32496B49998F247;
precomp_x[27] = 256'hCAF754272DC84563B0352B7A14311AF55D245315ACE27C65369E15F7151D41D1;
precomp_x[28] = 256'h2600CA4B282CB986F85D0F1709979D8B44A09C07CB86D7C124497BC86F082120;
precomp_x[29] = 256'h7635CA72D7E8432C338EC53CD12220BC01C48685E24F7DC8C602A7746998E435;
precomp_x[30] = 256'h754E3239F325570CDBBF4A87DEEE8A66B7F2B33479D468FBC1A50743BF56CC18;
precomp_x[31] = 256'hE3E6BD1071A1E96AFF57859C82D570F0330800661D1C952F9FE2694691D9B9E8;
precomp_y[0] = 256'h483ADA7726A3C4655DA4FBFC0E1108A8FD17B448A68554199C47D08FFB10D4B8;
precomp_y[1] = 256'h388F7B0F632DE8140FE337E62A37F3566500A99934C2231B6CB9FD7584B8E672;
precomp_y[2] = 256'hD8AC222636E5E3D6D4DBA9DDA6C9C426F788271BAB0D6840DCA87D3AA6AC62D6;
precomp_y[3] = 256'h6AEBCA40BA255960A3178D6D861A54DBA813D0B813FDE7B5A5082628087264DA;
precomp_y[4] = 256'hCC338921B0A7D9FD64380971763B61E9ADD888A4375F8E0F05CC262AC64F9C37;
precomp_y[5] = 256'hD984A032EB6B5E190243DD56D7B7B365372DB1E2DFF9D6A8301D74C9C953C61B;
precomp_y[6] = 256'h0AB0902E8D880A89758212EB65CDAF473A1A06DA521FA91F29B5CB52DB03ED81;
precomp_y[7] = 256'h581E2872A86C72A683842EC228CC6DEFEA40AF2BD896D3A5C504DC9FF6A26B58;
precomp_y[8] = 256'h4211AB0694635168E997B0EAD2A93DAECED1F4A04A95C0F6CFB199F69E56EB77;
precomp_y[9] = 256'h85E89BC037945D93B343083B5A1C86131A01F60C50269763B570C854E5C09B7A;
precomp_y[10] = 256'h321EB4075348F534D59C18259DDA3E1F4A1B3B2E71B1039C67BD3D8BCF81998C;
precomp_y[11] = 256'h02DE1068295DD865B64569335BD5DD80181D70ECFC882648423BA76B532B7D67;
precomp_y[12] = 256'h73016F7BF234AADE5D1AA71BDEA2B1FF3FC0DE2A887912FFE54A32CE97CB3402;
precomp_y[13] = 256'hA69DCE4A7D6C98E8D4A1ACA87EF8D7003F83C230F3AFA726AB40E52290BE1C55;
precomp_y[14] = 256'h2119A460CE326CDC76C45926C982FDAC0E106E861EDF61C5A039063F0E0E6482;
precomp_y[15] = 256'hE022CF42C2BD4A708B3F5126F16A24AD8B33BA48D0423B6EFD5E6348100D8A82;
precomp_y[16] = 256'hB9C398F186806F5D27561506E4557433A2CF15009E498AE7ADEE9D63D01B2396;
precomp_y[17] = 256'h02972D2DE4F8D20681A78D93EC96FE23C26BFAE84FB14DB43B01E1E9056B8C49;
precomp_y[18] = 256'h80FC06BD8CC5B01098088A1950EED0DB01AA132967AB472235F5642483B25EAF;
precomp_y[19] = 256'h1C38303F1CC5C30F26E66BAD7FE72F70A65EED4CBE7024EB1AA01F56430BD57A;
precomp_y[20] = 256'h0D0E3FA9ECA8726909559E0D79269046BDC59EA10C70CE2B02D499EC224DC7F7;
precomp_y[21] = 256'hEECF41253136E5F99966F21881FD656EBC4345405C520DBC063465B521409933;
precomp_y[22] = 256'h758F3F41AFD6ED428B3081B0512FD62A54C3F3AFBB5B6764B653052A12949C9A;
precomp_y[23] = 256'h958EF42A7886B6400A08266E9BA1B37896C95330D97077CBBE8EB3C7671C60D6;
precomp_y[24] = 256'hE0DEDC9B3B2F8DAD4DA1F32DEC2531DF9EB5FBEB0598E4FD1A117DBA703A3C37;
precomp_y[25] = 256'h5ED430D78C296C3543114306DD8622D7C622E27C970A1DE31CB377B01AF7307E;
precomp_y[26] = 256'hCEDABD9B82203F7E13D206FCDF4E33D92A6C53C26E5CCE26D6579962C4E31DF6;
precomp_y[27] = 256'hCB474660EF35F5F2A41B643FA5E460575F4FA9B7962232A5C32F908318A04476;
precomp_y[28] = 256'h4119B88753C15BD6A693B03FCDDBB45D5AC6BE74AB5F0EF44B0BE9475A7E4B40;
precomp_y[29] = 256'h091B649609489D613D1D5E590F78E6D74ECFC061D57048BAD9E76F302C5B9C61;
precomp_y[30] = 256'h0673FB86E5BDA30FB3CD0ED304EA49A023EE33D0197A695D0C5D98093C536683;
precomp_y[31] = 256'h59C9E0BBA394E76F40C0AA58379A3CB6A5A2283993E90C4167002AF4920E37F5;
