precomp_y[0] = 256'h483ADA7726A3C4655DA4FBFC0E1108A8FD17B448A68554199C47D08FFB10D4B8;
precomp_y[1] = 256'h388F7B0F632DE8140FE337E62A37F3566500A99934C2231B6CB9FD7584B8E672;
precomp_y[2] = 256'hD8AC222636E5E3D6D4DBA9DDA6C9C426F788271BAB0D6840DCA87D3AA6AC62D6;
precomp_y[3] = 256'h6AEBCA40BA255960A3178D6D861A54DBA813D0B813FDE7B5A5082628087264DA;
precomp_y[4] = 256'hCC338921B0A7D9FD64380971763B61E9ADD888A4375F8E0F05CC262AC64F9C37;
precomp_y[5] = 256'hD984A032EB6B5E190243DD56D7B7B365372DB1E2DFF9D6A8301D74C9C953C61B;
precomp_y[6] = 256'h0AB0902E8D880A89758212EB65CDAF473A1A06DA521FA91F29B5CB52DB03ED81;
precomp_y[7] = 256'h581E2872A86C72A683842EC228CC6DEFEA40AF2BD896D3A5C504DC9FF6A26B58;
precomp_y[8] = 256'h4211AB0694635168E997B0EAD2A93DAECED1F4A04A95C0F6CFB199F69E56EB77;
precomp_y[9] = 256'h85E89BC037945D93B343083B5A1C86131A01F60C50269763B570C854E5C09B7A;
precomp_y[10] = 256'h321EB4075348F534D59C18259DDA3E1F4A1B3B2E71B1039C67BD3D8BCF81998C;
precomp_y[11] = 256'h02DE1068295DD865B64569335BD5DD80181D70ECFC882648423BA76B532B7D67;
precomp_y[12] = 256'h73016F7BF234AADE5D1AA71BDEA2B1FF3FC0DE2A887912FFE54A32CE97CB3402;
precomp_y[13] = 256'hA69DCE4A7D6C98E8D4A1ACA87EF8D7003F83C230F3AFA726AB40E52290BE1C55;
precomp_y[14] = 256'h2119A460CE326CDC76C45926C982FDAC0E106E861EDF61C5A039063F0E0E6482;
precomp_y[15] = 256'hE022CF42C2BD4A708B3F5126F16A24AD8B33BA48D0423B6EFD5E6348100D8A82;
precomp_y[16] = 256'hB9C398F186806F5D27561506E4557433A2CF15009E498AE7ADEE9D63D01B2396;
precomp_y[17] = 256'h02972D2DE4F8D20681A78D93EC96FE23C26BFAE84FB14DB43B01E1E9056B8C49;
precomp_y[18] = 256'h80FC06BD8CC5B01098088A1950EED0DB01AA132967AB472235F5642483B25EAF;
precomp_y[19] = 256'h1C38303F1CC5C30F26E66BAD7FE72F70A65EED4CBE7024EB1AA01F56430BD57A;
precomp_y[20] = 256'h0D0E3FA9ECA8726909559E0D79269046BDC59EA10C70CE2B02D499EC224DC7F7;
precomp_y[21] = 256'hEECF41253136E5F99966F21881FD656EBC4345405C520DBC063465B521409933;
precomp_y[22] = 256'h758F3F41AFD6ED428B3081B0512FD62A54C3F3AFBB5B6764B653052A12949C9A;
precomp_y[23] = 256'h958EF42A7886B6400A08266E9BA1B37896C95330D97077CBBE8EB3C7671C60D6;
precomp_y[24] = 256'hE0DEDC9B3B2F8DAD4DA1F32DEC2531DF9EB5FBEB0598E4FD1A117DBA703A3C37;
precomp_y[25] = 256'h5ED430D78C296C3543114306DD8622D7C622E27C970A1DE31CB377B01AF7307E;
precomp_y[26] = 256'hCEDABD9B82203F7E13D206FCDF4E33D92A6C53C26E5CCE26D6579962C4E31DF6;
precomp_y[27] = 256'hCB474660EF35F5F2A41B643FA5E460575F4FA9B7962232A5C32F908318A04476;
precomp_y[28] = 256'h4119B88753C15BD6A693B03FCDDBB45D5AC6BE74AB5F0EF44B0BE9475A7E4B40;
precomp_y[29] = 256'h091B649609489D613D1D5E590F78E6D74ECFC061D57048BAD9E76F302C5B9C61;
precomp_y[30] = 256'h0673FB86E5BDA30FB3CD0ED304EA49A023EE33D0197A695D0C5D98093C536683;
precomp_y[31] = 256'h59C9E0BBA394E76F40C0AA58379A3CB6A5A2283993E90C4167002AF4920E37F5;
precomp_y[32] = 256'h3B952D32C67CF77E2E17446E204180AB21FB8090895138B4A4A797F86E80888B;
precomp_y[33] = 256'h55EB2DAFD84D6CCD5F862B785DC39D4AB157222720EF9DA217B8C45CF2BA2417;
precomp_y[34] = 256'hEFAE9C8DBC14130661E8CEC030C89AD0C13C66C0D17A2905CDC706AB7399A868;
precomp_y[35] = 256'hE38DA76DCD440621988D00BCF79AF25D5B29C094DB2A23146D003AFD41943E7A;
precomp_y[36] = 256'hF98A3FD831EB2B749A93B0E6F35CFB40C8CD5AA667A15581BC2FEDED498FD9C6;
precomp_y[37] = 256'h744B1152EACBE5E38DCC887980DA38B897584A65FA06CEDD2C924F97CBAC5996;
precomp_y[38] = 256'hC534AD44175FBC300F4EA6CE648309A042CE739A7919798CD85E216C4A307F6E;
precomp_y[39] = 256'hE13817B44EE14DE663BF4BC808341F326949E21A6A75C2570778419BDAF5733D;
precomp_y[40] = 256'h30E93E864E669D82224B967C3020B8FA8D1E4E350B6CBCC537A48B57841163A2;
precomp_y[41] = 256'hE491A42537F6E597D5D28A3224B1BC25DF9154EFBD2EF1D2CBBA2CAE5347D57E;
precomp_y[42] = 256'h100B610EC4FFB4760D5C1FC133EF6F6B12507A051F04AC5760AFA5B29DB83437;
precomp_y[43] = 256'hEF0AFBB2056205448E1652C48E8127FC6039E77C15C2378B7E7D15A0DE293311;
precomp_y[44] = 256'h8B378A22D827278D89C5E9BE8F9508AE3C2AD46290358630AFB34DB04EEDE0A4;
precomp_y[45] = 256'h68651CF9B6DA903E0914448C6CD9D4CA896878F5282BE4C8CC06E2A404078575;
precomp_y[46] = 256'hF5435A2BD2BADF7D485A4D8B8DB9FCCE3E1EF8E0201E4578C54673BC1DC5EA1D;
precomp_y[47] = 256'hD56EB30B69463E7234F5137B73B84177434800BACEBFC685FC37BBE9EFE4070D;
precomp_y[48] = 256'hEDD77F50BCB5A3CAB2E90737309667F2641462A54070F3D519212D39C197A629;
precomp_y[49] = 256'h0A855BABAD5CD60C88B430A69F53A1A7A38289154964799BE43D06D77D31DA06;
precomp_y[50] = 256'h66DB656F87D1F04FFFD1F04788C06830871EC5A64FEEE685BD80F0B1286D8374;
precomp_y[51] = 256'h09414685E97B1B5954BD46F730174136D57F1CEEB487443DC5321857BA73ABEE;
precomp_y[52] = 256'h4CB95957E83D40B0F73AF4544CCCF6B1F4B08D3C07B27FB8D8C2962A400766D1;
precomp_y[53] = 256'hFA77968128D9C92EE1010F337AD4717EFF15DB5ED3C049B3411E0315EAA4593B;
precomp_y[54] = 256'h5F3032F5892156E39CCD3D7915B9E1DA2E6DAC9E6F26E961118D14B8462E1661;
precomp_y[55] = 256'h8EC0BA238B96BEC0CBDDDCAE0AA442542EEE1FF50C986EA6B39847B3CC092FF6;
precomp_y[56] = 256'h8DC2412AAFE3BE5C4C5F37E0ECC5F9F6A446989AF04C4E25EBAAC479EC1C8C1E;
precomp_y[57] = 256'h5E4631150E62FB40D0E8C2A7CA5804A39D58186A50E497139626778E25B0674D;
precomp_y[58] = 256'hF65F5D3E292C2E0819A528391C994624D784869D7E6EA67FB18041024EDC07DC;
precomp_y[59] = 256'hF3E0319169EB9B85D5404795539A5E68FA1FBD583C064D2462B675F194A3DDB4;
precomp_y[60] = 256'h42242A969283A5F339BA7F075E36BA2AF925CE30D767ED6E55F4B031880D562C;
precomp_y[61] = 256'h204B5D6F84822C307E4B4A7140737AEC23FC63B65B35F86A10026DBD2D864E6B;
precomp_y[62] = 256'h04F14351D0087EFA49D245B328984989D5CAF9450F34BFC0ED16E96B58FA9913;
precomp_y[63] = 256'h073867F59C0659E81904F9A1C7543698E62562D6744C169CE7A36DE01A8D6154;
precomp_y[64] = 256'h39F23F366809085BEEBFC71181313775A99C9AED7D8BA38B161384C746012865;
precomp_y[65] = 256'hD2424B1B1ABE4EB8164227B085C9AA9456EA13493FD563E06FD51CF5694C78FC;
precomp_y[66] = 256'hEAD12168595FE1BE99252129B6E56B3391F7AB1410CD1E0EF3DCDCABD2FDA224;
precomp_y[67] = 256'h6FDCEF09F2F6D0A044E654AEF624136F503D459C3E89845858A47A9129CDD24E;
precomp_y[68] = 256'h060660257DD11B3AA9C8ED618D24EDFF2306D320F1D03010E33A7D2057F3B3B6;
precomp_y[69] = 256'h3D98A9CDD026DD43F39048F25A8847F4FCAFAD1895D7A633C6FED3C35E999511;
precomp_y[70] = 256'h0B4C4FE99C775A606E2D8862179139FFDA61DC861C019E55CD2876EB2A27D84B;
precomp_y[71] = 256'hAE434102EDDE0958EC4B19D917A6A28E6B72DA1834AFF0E650F049503A296CF2;
precomp_y[72] = 256'hCF2174118C8B6D7A4B48F6D534CE5C79422C086A63460502B827CE62A326683C;
precomp_y[73] = 256'h6FB8D5591B466F8FC63DB50F1C0F1C69013F996887B8244D2CDEC417AFEA8FA3;
precomp_y[74] = 256'h322AF4908C7312B0CFBFE369F7A7B3CDB7D4494BC2823700CFD652188A3EA98D;
precomp_y[75] = 256'h6749E67C029B85F52A034EAFD096836B2520818680E26AC8F3DFBCDB71749700;
precomp_y[76] = 256'h2AEABE7E4531510116217F07BF4D07300DE97E4874F81F533420A72EEB0BD6A4;
precomp_y[77] = 256'hB0EA558A113C30BEA60FC4775460C7901FF0B053D25CA2BDEEE98F1A4BE5D196;
precomp_y[78] = 256'h998C74A8CD45AC01289D5833A7BEB4744FF536B01B257BE4C5767BEA93EA57A4;
precomp_y[79] = 256'hB2284279995A34E2F9D4DE7396FC18B80F9B8B9FDD270F6661F79CA4C81BD257;
precomp_y[80] = 256'hBDD46039FEED17881D1E0862DB347F8CF395B74FC4BCDC4E940B74E3AC1F1B13;
precomp_y[81] = 256'h6F0A256BC5EFDF429A2FB6242F1A43A2D9B925BB4A4B3A26BB8E0F45EB596096;
precomp_y[82] = 256'hC359D6923BB398F7FD4473E16FE1C28475B740DD098075E6C0E8649113DC3A38;
precomp_y[83] = 256'h021AE7F4680E889BB130619E2C0F95A360CEB573C70603139862AFD617FA9B9F;
precomp_y[84] = 256'h60EA7F61A353524D1C987F6ECEC92F086D565AB687870CB12689FF1E31C74448;
precomp_y[85] = 256'h49B96715AB6878A79E78F07CE5680C5D6673051B4935BD897FEA824B77DC208A;
precomp_y[86] = 256'h5CA560753BE2A12FC6DE6CAF2CB489565DB936156B9514E1BB5E83037E0FA2D4;
precomp_y[87] = 256'h7571D74EE5E0FB92A7A8B33A07783341A5492144CC54BCC40A94473693606437;
precomp_y[88] = 256'hBE52D107BCFA09D8BCB9736A828CFA7FAC8DB17BF7A76A2C42AD961409018CF7;
precomp_y[89] = 256'h8FD64A14C06B589C26B947AE2BCF6BFA0149EF0BE14ED4D80F448A01C43B1C6D;
precomp_y[90] = 256'h39E5C9925B5A54B07433A4F18C61726F8BB131C012CA542EB24A8AC07200682A;
precomp_y[91] = 256'h62DFAF07A0F78FEB30E30D6295853CE189E127760AD6CF7FAE164E122A208D54;
precomp_y[92] = 256'h25A748AB367979D98733C38A1FA1C2E7DC6CC07DB2D60A9AE7A76AAA49BD0F77;
precomp_y[93] = 256'hECFB7056CF1DE042F9420BAB396793C0C390BDE74B4BBDFF16A83AE09A9A7517;
precomp_y[94] = 256'hCD450EC335438986DFEFA10C57FEA9BCC521A0959B2D80BBF74B190DCA712D10;
precomp_y[95] = 256'hF5C54754A8F71EE540B9B48728473E314F729AC5308B06938360990E2BFAD125;
precomp_y[96] = 256'h6CB9A8876D9CB8520609AF3ADD26CD20A0A7CD8A9411131CE85F44100099223E;
precomp_y[97] = 256'hFEF5A3C68059A6DEC5D624114BF1E91AAC2B9DA568D6ABEB2570D55646B8ADF1;
precomp_y[98] = 256'h1ACB250F255DD61C43D94CCC670D0F58F49AE3FA15B96623E5430DA0AD6C62B2;
precomp_y[99] = 256'h5F310D4B3C99B9EBB19F77D41C1DEE018CF0D34FD4191614003E945A1216E423;
precomp_y[100] = 256'h438136D603E858A3A5C440C38ECCBADDC1D2942114E2EDDD4740D098CED1F0D8;
precomp_y[101] = 256'hCDB559EEDC2D79F926BAF44FB84EA4D44BCF50FEE51D7CEB30E2E7F463036758;
precomp_y[102] = 256'h0C3B997D050EE5D423EBAF66A6DB9F57B3180C902875679DE924B69D84A7B375;
precomp_y[103] = 256'h6D89AD7BA4876B0B22C2CA280C682862F342C8591F1DAF5170E07BFD9CCAFA7D;
precomp_y[104] = 256'hCA5EF7D4B231C94C3B15389A5F6311E9DAFF7BB67B103E9880EF4BFF637ACAEC;
precomp_y[105] = 256'h09731141D81FC8F8084D37C6E7542006B3EE1B40D60DFE5362A5B132FD17DDC0;
precomp_y[106] = 256'hEE1849F513DF71E32EFC3896EE28260C73BB80547AE2275BA497237794C8753C;
precomp_y[107] = 256'hD3AA2ED71C9DD2247A62DF062736EB0BADDEA9E36122D2BE8641ABCB005CC4A4;
precomp_y[108] = 256'hC4E1020916980A4DA5D01AC5E6AD330734EF0D7906631C4F2390426B2EDD791F;
precomp_y[109] = 256'h67163E903236289F776F22C25FB8A3AFC1732F2B84B4E95DBDA47AE5A0852649;
precomp_y[110] = 256'h0CD1BC7CB6CC407BB2F0CA647C718A730CF71872E7D0D2A53FA20EFCDFE61826;
precomp_y[111] = 256'h299D21F9413F33B3EDF43B257004580B70DB57DA0B182259E09EECC69E0D38A5;
precomp_y[112] = 256'hF9429E738B8E53B968E99016C059707782E14F4535359D582FC416910B3EEA87;
precomp_y[113] = 256'h462F9BCE619898638499350113BBC9B10A878D35DA70740DC695A559EB88DB7B;
precomp_y[114] = 256'h62188BC49D61E5428573D48A74E1C655B1C61090905682A0D5558ED72DCCB9BC;
precomp_y[115] = 256'h7C10DFB164C3425F5C71A3F9D7992038F1065224F72BB9D1D902A6D13037B47C;
precomp_y[116] = 256'hAB8C1E086D04E813744A655B2DF8D5F83B3CDC6FAA3088C1D3AEA1454E3A1D5F;
precomp_y[117] = 256'h4CB04437F391ED73111A13CC1D4DD0DB1693465C2240480D8955E8592F27447A;
precomp_y[118] = 256'hBD1AEB21AD22EBB22A10F0303417C6D964F8CDD7DF0ACA614B10DC14D125AC46;
precomp_y[119] = 256'hBFEFACDB0E5D0FD7DF3A311A94DE062B26B80C61FBC97508B79992671EF7CA7F;
precomp_y[120] = 256'h603C12DAF3D9862EF2B25FE1DE289AED24ED291E0EC6708703A5BD567F32ED03;
precomp_y[121] = 256'hCC6157EF18C9C63CD6193D83631BBEA0093E0968942E8C33D5737FD790E0DB08;
precomp_y[122] = 256'h553E04F6B018B4FA6C8F39E7F311D3176290D0E0F19CA73F17714D9977A22FF8;
precomp_y[123] = 256'h0712FCDD1B9053F09003A3481FA7762E9FFD7C8EF35A38509E2FBF2629008373;
precomp_y[124] = 256'hED8CC9D04B29EB877D270B4878DC43C19AEFD31F4EEE09EE7B47834C1FA4B1C3;
precomp_y[125] = 256'h9852390A99507679FD0B86FD2B39A868D7EFC22151346E1A3CA4726586A6BED8;
precomp_y[126] = 256'h9E994980D9917E22B76B061927FA04143D096CCC54963E6A5EBFA5F3F8E286C1;
precomp_y[127] = 256'h4036EDC931A60AE889353F77FD53DE4A2708B26B6F5DA72AD3394119DAF408F9;
precomp_y[128] = 256'h753C8B9F9754F18D87F21145D9E2936B5EE050B27BBD9681442C76E92FCF91E6;
precomp_y[129] = 256'h86CA160D68F4D4E718B495B891D3B1B573B871A702B4CF6123ABD4483AA79C64;
precomp_y[130] = 256'h8147CBF7B973FCC15B57B6A3CFAD6863EDD0F30E3C45B85DC300C513C247759D;
precomp_y[131] = 256'h31B3CA455073BEA558ADBE56C27B470BAF949AE650213921DC287844F1A29574;
precomp_y[132] = 256'h57FC24472225B23F5714626D8D67D56110BD3A60DD7A16870CBBB893F652F50F;
precomp_y[133] = 256'h844ADB5CE7D10DE94617C73CA77040E4EE4E92E0156B3C70CC593FA494B33482;
precomp_y[134] = 256'hD765466C6E556E352F77872225627D80A73538074B44FF27057AD22E2F2454A2;
precomp_y[135] = 256'h77B1F0687CFCDBE8812605E50D8B752CDA811844236A4C4377F53C946E7BD648;
precomp_y[136] = 256'hC16F60C7C11FC3C9EB27FA26A9035B669BFB77D21CEF371DDCE94E329222550C;
precomp_y[137] = 256'hE1BCFE7FC8ED8AE95CF6C2437FDD94BFD742E8CAA6DE78114C25112A86988EFD;
precomp_y[138] = 256'h8D6857C9D08EF7B4FD8883363D37BEE70FE8529F7173F58943FCAE81D2D0EA0E;
precomp_y[139] = 256'hDDF1B9FE8744AD03F996BF6B96EC34962B601BD5ED952F7854F583888917BE80;
precomp_y[140] = 256'h3F27E7E1834F1A61AF6F04DC61E7AE64716BC5E0A6B063B301D0E60E47298A9D;
precomp_y[141] = 256'h50BC23F3926CD0C49F53FBB235EB1E890D579517F5BDC3AB2416DB785AAEDB3F;
precomp_y[142] = 256'h6E6AEE6C9625370AF866C25C7CA5DD780527EFBCE7D8B3A39AB249309A185187;
precomp_y[143] = 256'h986314EF75B68FB2827C2965041981395D699FCD81CF23CE7019BC4135174870;
precomp_y[144] = 256'h4E31EA12AC607D075DE4B22DE1BE2C52E0A44D254728D2C544D2DDF9E3E469C0;
precomp_y[145] = 256'h94264621A5960E0EE24C27926F16CAD2907F2636762E8D5A17E94AFD8E9D2BB0;
precomp_y[146] = 256'h5B5853AB7EE5DE8D34E3D6BEB201094FFF8FBD1E0682F7F1EF87DDD65D7303C9;
precomp_y[147] = 256'h496C944DD9875BA60A537EF96BF4C714A0AFFF24387D95E89B42337A33110753;
precomp_y[148] = 256'hF2ECCAC775922B50899C979A02B3CC30B629E62E85693BA470F6EE381284C162;
precomp_y[149] = 256'h44C757A542F4EA2EB39605D4268C2510AC685AABD77A8F5C4D95E23F4C2E9368;
precomp_y[150] = 256'h7421A2207EE73299D46192FC93CA03DEC824ED8DE2F48367EC5383170A17FFFB;
precomp_y[151] = 256'h7D16D654F0C2AFF0FC254DAD063761A26C8D4022EA85B8CC22F3EA1EF69961A9;
precomp_y[152] = 256'h6C9ED1F1528B021593A39839340DDB530A2F2E365290C49824B035C673C9259D;
precomp_y[153] = 256'h0E8BCBFE1F7F6E75D32E20499329765F02EFFC56A922F26860D4BC0AADD0E24D;
precomp_y[154] = 256'h3E18941CC3C6D297CC9A32F695807B1C7DA8561DE4FDE71D4F9BBDB6E9BF3916;
precomp_y[155] = 256'hF60547AB6E9C5FD3ECA6E349B85880C61FDAD0FC2F7AB155295CAAECB973C154;
precomp_y[156] = 256'h29A835F6EF7FA1E5F6F37A80CF96CA9843762BB1B12A0DAEAE83234BD0B5CCD5;
precomp_y[157] = 256'h5C7BCF8B57F114E0B73BCFB810F5C60D35DC99AE9DC7F0E2606CC1F728C2071E;
precomp_y[158] = 256'hA286E222DFE10CFD9689EABA6A81F04489C86DB6869AA1B554A90F1E83778EEE;
precomp_y[159] = 256'hC582DB1A3F0F22421913B2E951E98A78660B4C40AD08FD65528593BC18223188;
precomp_y[160] = 256'hE3E77C41288F2602E722AF7F4B70E64DE4116FB9955B03B06EA8B19F7A20350D;
precomp_y[161] = 256'hC9E33FAEBD8EBA426736C0C76F3DEABAEE2B59C50953FB43C2DCC5139E7C4BDC;
precomp_y[162] = 256'hF5202CF5AAEEA58BF4F58C7EDF4417BE1B87FFDEE68E77F0D7E81ABE158E3A25;
precomp_y[163] = 256'h61FE64CAB0952CAE3C574F282F74A87DC2A96316B7009F2E4E9C5FCC12285844;
precomp_y[164] = 256'h5DCF9ABBA9625ED680B0F20FB1F047D593A0C61C539692538CDF6B034D730B58;
precomp_y[165] = 256'h79A6BF4375F1469C4F5321C6C72FBBF4BA7CEC105675F437B5E013AD7B5D75D4;
precomp_y[166] = 256'h7669BBD419A4D491F592A35B6AA3DFE45BD2FE7FD179C7781CD5F918D732F63D;
precomp_y[167] = 256'h308ABC8DF271F75959B20C5C7FA62BAFBFC9CCBF49B946A954E5381C1728D1C7;
precomp_y[168] = 256'h9EEA970BA856B2FAA3E82877CC84ED4F3DC0EFBA1E7C3BAA8B386FFC46E0AE7E;
precomp_y[169] = 256'hA9FB1702100953B359B2E2688AE7FD33A30377DA47BFDA713E2D7D73DFB1030C;
precomp_y[170] = 256'h22F6FE9D217495017FDB7F5B2F12FA57095F40E131714885C12A2EA16EDB6BE6;
precomp_y[171] = 256'h737CECA2C0EF72278B90501CCB71B6715E5C31D4CD0478C118FE128795F1DD0C;
precomp_y[172] = 256'h2AFC8D09B79176D8D003FD2A4F18D526403FFF272D47E7787376FEB7CBDDD8FD;
precomp_y[173] = 256'hCB13C152FD511D91A9E0ED90AFA021A081F77F6D20CC1376E2195FFCF28FA758;
precomp_y[174] = 256'h1AB4EABE5E09409D75CCA8922647F48DBD698A16D4F7CC8596DAF16940023A52;
precomp_y[175] = 256'h95F9F4E9007E5B9FA48FA422A26AB982DC48A4D54D7123986E6D3AB974E88915;
precomp_y[176] = 256'hDCE1BAE1D655BA517F5B5580997117570A77CD3BDD4B8E8E330E97791BC31DF0;
precomp_y[177] = 256'hCC3636A03FDDDDFABED88DAAB081F3591C48D2CA71BA34FCF6989F4AF7625D8E;
precomp_y[178] = 256'h329CF0497E15EEC7B8EAFC4A0B8A7D1CD8B632038D4AEF81974CF9844611A32D;
precomp_y[179] = 256'h8C6F81BE3FAFA5EEC8296F928AC7919DC4D88C9A59442274D0531B7BF7E48E78;
precomp_y[180] = 256'h7F42C0962FEB2F73B2B0965A1F359A6ADE49D768A2CE6B07B5ACB92B73E05583;
precomp_y[181] = 256'hF649BE278CAD976420742CE382DCE3A1420E372EF1B25B2759A8ED387282765E;
precomp_y[182] = 256'hD596ADF0E8692A06BC6284BF0299BEF685E2A171585AA1324B9A05B50CE815B7;
precomp_y[183] = 256'hE077184B4AE8F7056C10DD9EF541689D143F6871789E1801DEAEFC1D527A8FB4;
precomp_y[184] = 256'hEB4C98489093D573A295407E1D6FC48A787120CEB3D3DCFBB40634E0E75E221D;
precomp_y[185] = 256'hEA75B9B25D717861D1AF1C019C372941C8968B90EF134F9F323215E1BB0B2155;
precomp_y[186] = 256'h669985206EDF4AC6F39BE21F20C98824210E204CE44998095DE355371641218C;
precomp_y[187] = 256'h70B0123774AF550E68E68E5F65CA6E9808846E03CF39AF778511BE82BC32FEFE;
precomp_y[188] = 256'hE115B14BEF4695CFFB85BDF98BA3985CBD5E5B8983E053907C36F9CE8B75D41D;
precomp_y[189] = 256'hE9D9DBFE8CF5F5CCA855D6CCBD11F48060FAFA8DAD6BD3E9C86DF5CEB0FA5270;
precomp_y[190] = 256'hE4177CE1C3CD6AC778925BD67E72CB77D1925B91D06A7F1698411A4786393FB0;
precomp_y[191] = 256'h954A5FD857BA3ACF2D4B1F41E8E1F2CD1F21C4B96899781B742A49D2E61ED18B;
precomp_y[192] = 256'h2D5D2FB1F0C308553B1FE249298B2059259D3D49D4D7071ADCE4BCC5DC937193;
precomp_y[193] = 256'h9BD0178E381895692217267B7407E98727FCAEDA12D8CF5449EB5472D554E0FF;
precomp_y[194] = 256'h618BD6B0D25CA70DF08B76929336E421691B09730F2F5A052E7ADC173584427B;
precomp_y[195] = 256'h07A981F0C21862A853B4F895DC62482C530ED7385E5D1E330CFB9D0FE879992C;
precomp_y[196] = 256'hADB23BCDB3D069C5E83BE30B2469B0680B2A81B7B667E934233B75EFB5753F28;
precomp_y[197] = 256'hD8003C9EE3C842F5EDE375A8A7768DB4803ECF119B7B37DECEA15631B4E8DBCA;
precomp_y[198] = 256'h211557489FA93B883E5BEA50DA005C5368E21A0C41BC83D9145C13E1370D26D0;
precomp_y[199] = 256'hABB1D9F874637668E214EFBAFBF529D312FF023BC1D5723E585404366834F189;
precomp_y[200] = 256'h5B5930F12E9C40BCB3393A895C2D64576A3ABD23B7291B99C965C33DEF60A55C;
precomp_y[201] = 256'h5246A8190BBFB2915F82ED5650796F505CED5C2587347D57A873CEAF3D997E7A;
precomp_y[202] = 256'h3C83145DAD9F87487B97E7464850ED02D71DBD04093281A13D2127766A791EE2;
precomp_y[203] = 256'h6CE693B64A37C6727E141041AB9A0D589AB9C303A5AC3D3EC89B6F279E79827C;
precomp_y[204] = 256'hF602C3428593A9A8D671D1BC7C1D88340FE9F5F52E6A7F0FBB8701464E6F4838;
precomp_y[205] = 256'hB8F7C3B220701320F20CA036761D3E56BF94A7009A919F1A3EA0CB81B74424A6;
precomp_y[206] = 256'hAFB6A74D9849454EDD7F703A5C6616D143F9CBCC9A9A5D6F6A7B5D1F9D9FCAFF;
precomp_y[207] = 256'hDA7D67CBC1EDE9D4FEDD5DCDC96B04F9A3561BA02581B055EAA144EB4217DACA;
precomp_y[208] = 256'h160E1C1C13342FD459D4F9898AE632B842B8947913733B89384FC1042D30BF01;
precomp_y[209] = 256'h87092DCBB9C3D254E3B055FF3A76EC0564C4A7C57FB1783CEFDC40FC10B751F0;
precomp_y[210] = 256'hFE49A6A8B5E46BF1EF679714DABD590EA831D46B8EE94EB613132BA37855FABB;
precomp_y[211] = 256'h4521954EFCC98263DF2F14E0E6E6B47AF6B83F0BBC20722C15445F87E05F4513;
precomp_y[212] = 256'hCD15ABBCD744D4850D5E401F1F89A5DF122F37B4E362B4CEE3E53B1C00110BF3;
precomp_y[213] = 256'hCFD4D36BEB2E11F241FD0F367A0737AD303E915FF247F131368CA50918E00957;
precomp_y[214] = 256'h72EA16B532A7336D3332400B303C0236B6A1294D88CE7FE915571284D1F7C189;
precomp_y[215] = 256'hD5E6268B30952422BE59FE0EFE7BA2E703215994827A46C2F2972B26153CF7AE;
precomp_y[216] = 256'hB8241453ABC44C57DDAD6FF386D416F43E258A390C6F88379F80472B943F32B9;
precomp_y[217] = 256'hC1FDAC5AEF4C6F0FFCB8E1C5C4417C713E3D5F07146DAA1AAAF2E7FEE70C4914;
precomp_y[218] = 256'hFD5A31976FAD6AEEC304752CC3EBBC511F3695B09A737FA30AF42CC6EFD684CC;
precomp_y[219] = 256'h563651760897632F8DDE31677A24F55834C5C9A55C1CBF36FD8B44803C9C6C81;
precomp_y[220] = 256'hB5CE31605D6DD9C622CAE425CCD28912C4439820C06950CD4C86D9B453ABD7ED;
precomp_y[221] = 256'h933D348378A71F443788194AAFC545E7F53E37A6F779F96E8FA14CCDEDE3B4EB;
precomp_y[222] = 256'h2A7D3701A8724B12BD7C4830224AC083CBEA83D0543B541480BA8C8AE7731232;
precomp_y[223] = 256'hEA90F8AAE214EE16ED608A72366998994E311DC7780EF885B29290C3823C470E;
precomp_y[224] = 256'hCB7571C4071C552765BD289EA3CF3F38796DA2B12C953D0B8705125C4861D598;
precomp_y[225] = 256'h7BBBB198EB39973B76D87F8194D45150A66D4F3B128A40BEC989A405AD7C287B;
precomp_y[226] = 256'hA2F2F02A8272DE6E3DC8B39508959AD251B6D3D004C8195259A501E28FF7892A;
precomp_y[227] = 256'h8613BB848398681D66F1E75D5B6EF44FD827B6290F4956A441D8F503DD32B289;
precomp_y[228] = 256'h838E779334AA6FE6CAE90A62D359C339187B403215D97CDA4E62724AA5A50306;
precomp_y[229] = 256'h01FCABF21E19CE68EE12A3D284BD1304010FA5F5D45F9C15D4070243A8433047;
precomp_y[230] = 256'hE15723EB0E0BDBE6D6F28D6DA0443C634851F5B4C551BEC69F9196A00969ED71;
precomp_y[231] = 256'hFFB0E211C79FBB7978BD4E53A05A267FF1E32C34D6287DEE64576D31AB959AB2;
precomp_y[232] = 256'hF6A9186FF147B9B5FFC844B2EC0E255A1AE5537D75624288CE8421F87E94E1A4;
precomp_y[233] = 256'h8791C0007C09C94DB328034B88C5BBBC113335366679EB099A5E75B583BC2C2A;
precomp_y[234] = 256'h4B985B13C54990267FF564D2D4649C6F7E8FDBE1BA101D941C034E1464877B20;
precomp_y[235] = 256'h31CE61A87834F52EFCF8703F93696F425813015563CA5D9CE92D8FC281135B0D;
precomp_y[236] = 256'hBEA2A060505C13BC317CA083C5A8B85C9EAD5F6E1AC23FBEAC7CECEA9251C791;
precomp_y[237] = 256'h74962C3FED9A6E9C896635EA855323B608850091F84DEE333CDFF8D0D2827928;
precomp_y[238] = 256'h1CBCF83EA363E0D93E6ECC328653BA7AA165C526765B09F0696B0D61F122DB3A;
precomp_y[239] = 256'hD10B5A637AB546BFCC610E2D1C3D61F461B0A806E7BA29C73D3DE909E9FAE659;
precomp_y[240] = 256'h7B148EF273E1B131341AD4779342C7BC7B945A2CB52C448E4BB5FD503CEA1A19;
precomp_y[241] = 256'h5847F4E06C6530335E29EA94389EE3E6D916314A60126028650AB9E0BFCFBBA7;
precomp_y[242] = 256'h2CBFAD4D16C0702186611EEC408082FBFB2E9898141A52481C59E44ECD0676FF;
precomp_y[243] = 256'h328E831D2F2B162C4ABE1644BB54CC8518DB178C5B6AE97E5E85110C7D7FDF1D;
precomp_y[244] = 256'h627EEA93C6C9B53F9455941440A8B1006EBA68D46C922B6A1521F3946DD15E4E;
precomp_y[245] = 256'h195A6A65D3790BEC716429863BCEF432E38242FC9F565DBBE159BC42F5740C69;
precomp_y[246] = 256'h177C3A61682363ABBF281615D59F06FF5F87644C84D670E9A6C56AC1B611509B;
precomp_y[247] = 256'h2D1A0B9C8EABA06543204DF148EB161825443EFA80F8AFF3D49B6626C5955AC8;
precomp_y[248] = 256'h549B18C310FEAEA10225FADE934112D34058101D74F005381B82796AD0461736;
precomp_y[249] = 256'hE95E050881AF550D09221F5AE95410316367D24BD545BDCB434E7638ACB46DBD;
precomp_y[250] = 256'h62F637C67D8863748F1E2E26865118B999285B8755F25512C968B4FE49B8C971;
precomp_y[251] = 256'hA0CBC0165E32171C8184265EAC7E0147206349D541035A94F56EFC49DCD7AB93;
precomp_y[252] = 256'hA532D00D35013F859F4041D3AA231F2B9FC499670E0E2F824D5051F9E7F0C626;
precomp_y[253] = 256'h92C20846CFDF1E8F3FE5BCAA06BDEDC39926833A3F40D28F23A8F952D8D18DDE;
precomp_y[254] = 256'h1F023F2FA2BBECE703DBA14C124095CBFDC4F92F00281A148304A412C16ECAE6;
precomp_y[255] = 256'h2DC6CAE5CAC2D88783DCA0E503C798F8FE067BCF5FC2975113756CF7EF4E5F1B;
precomp_x[0] = 256'h79BE667EF9DCBBAC55A06295CE870B07029BFCDB2DCE28D959F2815B16F81798;
precomp_x[1] = 256'hF9308A019258C31049344F85F89D5229B531C845836F99B08601F113BCE036F9;
precomp_x[2] = 256'h2F8BDE4D1A07209355B4A7250A5C5128E88B84BDDC619AB7CBA8D569B240EFE4;
precomp_x[3] = 256'h5CBDF0646E5DB4EAA398F365F2EA7A0E3D419B7E0330E39CE92BDDEDCAC4F9BC;
precomp_x[4] = 256'hACD484E2F0C7F65309AD178A9F559ABDE09796974C57E714C35F110DFC27CCBE;
precomp_x[5] = 256'h774AE7F858A9411E5EF4246B70C65AAC5649980BE5C17891BBEC17895DA008CB;
precomp_x[6] = 256'hF28773C2D975288BC7D1D205C3748651B075FBC6610E58CDDEEDDF8F19405AA8;
precomp_x[7] = 256'hD7924D4F7D43EA965A465AE3095FF41131E5946F3C85F79E44ADBCF8E27E080E;
precomp_x[8] = 256'hDEFDEA4CDB677750A420FEE807EACF21EB9898AE79B9768766E4FAA04A2D4A34;
precomp_x[9] = 256'h2B4EA0A797A443D293EF5CFF444F4979F06ACFEBD7E86D277475656138385B6C;
precomp_x[10] = 256'h352BBF4A4CDD12564F93FA332CE333301D9AD40271F8107181340AEF25BE59D5;
precomp_x[11] = 256'h2FA2104D6B38D11B0230010559879124E42AB8DFEFF5FF29DC9CDADD4ECACC3F;
precomp_x[12] = 256'h9248279B09B4D68DAB21A9B066EDDA83263C3D84E09572E269CA0CD7F5453714;
precomp_x[13] = 256'hDAED4F2BE3A8BF278E70132FB0BEB7522F570E144BF615C07E996D443DEE8729;
precomp_x[14] = 256'hC44D12C7065D812E8ACF28D7CBB19F9011ECD9E9FDF281B0E6A3B5E87D22E7DB;
precomp_x[15] = 256'h6A245BF6DC698504C89A20CFDED60853152B695336C28063B61C65CBD269E6B4;
precomp_x[16] = 256'h1697FFA6FD9DE627C077E3D2FE541084CE13300B0BEC1146F95AE57F0D0BD6A5;
precomp_x[17] = 256'h605BDB019981718B986D0F07E834CB0D9DEB8360FFB7F61DF982345EF27A7479;
precomp_x[18] = 256'h62D14DAB4150BF497402FDC45A215E10DCB01C354959B10CFE31C7E9D87FF33D;
precomp_x[19] = 256'h80C60AD0040F27DADE5B4B06C408E56B2C50E9F56B9B8B425E555C2F86308B6F;
precomp_x[20] = 256'h7A9375AD6167AD54AA74C6348CC54D344CC5DC9487D847049D5EABB0FA03C8FB;
precomp_x[21] = 256'hD528ECD9B696B54C907A9ED045447A79BB408EC39B68DF504BB51F459BC3FFC9;
precomp_x[22] = 256'h049370A4B5F43412EA25F514E8ECDAD05266115E4A7ECB1387231808F8B45963;
precomp_x[23] = 256'h77F230936EE88CBBD73DF930D64702EF881D811E0E1498E2F1C13EB1FC345D74;
precomp_x[24] = 256'hF2DAC991CC4CE4B9EA44887E5C7C0BCE58C80074AB9D4DBAEB28531B7739F530;
precomp_x[25] = 256'h463B3D9F662621FB1B4BE8FBBE2520125A216CDFC9DAE3DEBCBA4850C690D45B;
precomp_x[26] = 256'hF16F804244E46E2A09232D4AFF3B59976B98FAC14328A2D1A32496B49998F247;
precomp_x[27] = 256'hCAF754272DC84563B0352B7A14311AF55D245315ACE27C65369E15F7151D41D1;
precomp_x[28] = 256'h2600CA4B282CB986F85D0F1709979D8B44A09C07CB86D7C124497BC86F082120;
precomp_x[29] = 256'h7635CA72D7E8432C338EC53CD12220BC01C48685E24F7DC8C602A7746998E435;
precomp_x[30] = 256'h754E3239F325570CDBBF4A87DEEE8A66B7F2B33479D468FBC1A50743BF56CC18;
precomp_x[31] = 256'hE3E6BD1071A1E96AFF57859C82D570F0330800661D1C952F9FE2694691D9B9E8;
precomp_x[32] = 256'h186B483D056A033826AE73D88F732985C4CCB1F32BA35F4B4CC47FDCF04AA6EB;
precomp_x[33] = 256'hDF9D70A6B9876CE544C98561F4BE4F725442E6D2B737D9C91A8321724CE0963F;
precomp_x[34] = 256'h5EDD5CC23C51E87A497CA815D5DCE0F8AB52554F849ED8995DE64C5F34CE7143;
precomp_x[35] = 256'h290798C2B6476830DA12FE02287E9E777AA3FBA1C355B17A722D362F84614FBA;
precomp_x[36] = 256'hAF3C423A95D9F5B3054754EFA150AC39CD29552FE360257362DFDECEF4053B45;
precomp_x[37] = 256'h766DBB24D134E745CCCAA28C99BF274906BB66B26DCF98DF8D2FED50D884249A;
precomp_x[38] = 256'h59DBF46F8C94759BA21277C33784F41645F7B44F6C596A58CE92E666191ABE3E;
precomp_x[39] = 256'hF13ADA95103C4537305E691E74E9A4A8DD647E711A95E73CB62DC6018CFD87B8;
precomp_x[40] = 256'h7754B4FA0E8ACED06D4167A2C59CCA4CDA1869C06EBADFB6488550015A88522C;
precomp_x[41] = 256'h948DCADF5990E048AA3874D46ABEF9D701858F95DE8041D2A6828C99E2262519;
precomp_x[42] = 256'h7962414450C76C1689C7B48F8202EC37FB224CF5AC0BFA1570328A8A3D7C77AB;
precomp_x[43] = 256'h3514087834964B54B15B160644D915485A16977225B8847BB0DD085137EC47CA;
precomp_x[44] = 256'hD3CC30AD6B483E4BC79CE2C9DD8BC54993E947EB8DF787B442943D3F7B527EAF;
precomp_x[45] = 256'h1624D84780732860CE1C78FCBFEFE08B2B29823DB913F6493975BA0FF4847610;
precomp_x[46] = 256'h733CE80DA955A8A26902C95633E62A985192474B5AF207DA6DF7B4FD5FC61CD4;
precomp_x[47] = 256'h15D9441254945064CF1A1C33BBD3B49F8966C5092171E699EF258DFAB81C045C;
precomp_x[48] = 256'hA1D0FCF2EC9DE675B612136E5CE70D271C21417C9D2B8AAAAC138599D0717940;
precomp_x[49] = 256'hE22FBE15C0AF8CCC5780C0735F84DBE9A790BADEE8245C06C7CA37331CB36980;
precomp_x[50] = 256'h311091DD9860E8E20EE13473C1155F5F69635E394704EAA74009452246CFA9B3;
precomp_x[51] = 256'h34C1FD04D301BE89B31C0442D3E6AC24883928B45A9340781867D4232EC2DBDF;
precomp_x[52] = 256'hF219EA5D6B54701C1C14DE5B557EB42A8D13F3ABBCD08AFFCC2A5E6B049B8D63;
precomp_x[53] = 256'hD7B8740F74A8FBAAB1F683DB8F45DE26543A5490BCA627087236912469A0B448;
precomp_x[54] = 256'h32D31C222F8F6F0EF86F7C98D3A3335EAD5BCD32ABDD94289FE4D3091AA824BF;
precomp_x[55] = 256'h7461F371914AB32671045A155D9831EA8793D77CD59592C4340F86CBC18347B5;
precomp_x[56] = 256'hEE079ADB1DF1860074356A25AA38206A6D716B2C3E67453D287698BAD7B2B2D6;
precomp_x[57] = 256'h16EC93E447EC83F0467B18302EE620F7E65DE331874C9DC72BFD8616BA9DA6B5;
precomp_x[58] = 256'hEAA5F980C245F6F038978290AFA70B6BD8855897F98B6AA485B96065D537BD99;
precomp_x[59] = 256'h078C9407544AC132692EE1910A02439958AE04877151342EA96C4B6B35A49F51;
precomp_x[60] = 256'h494F4BE219A1A77016DCD838431AEA0001CDC8AE7A6FC688726578D9702857A5;
precomp_x[61] = 256'hA598A8030DA6D86C6BC7F2F5144EA549D28211EA58FAA70EBF4C1E665C1FE9B5;
precomp_x[62] = 256'hC41916365ABB2B5D09192F5F2DBEAFEC208F020F12570A184DBADC3E58595997;
precomp_x[63] = 256'h841D6063A586FA475A724604DA03BC5B92A2E0D2E0A36ACFE4C73A5514742881;
precomp_x[64] = 256'h5E95BB399A6971D376026947F89BDE2F282B33810928BE4DED112AC4D70E20D5;
precomp_x[65] = 256'h36E4641A53948FD476C39F8A99FD974E5EC07564B5315D8BF99471BCA0EF2F66;
precomp_x[66] = 256'h0336581EA7BFBBB290C191A2F507A41CF5643842170E914FAEAB27C2C579F726;
precomp_x[67] = 256'h8AB89816DADFD6B6A1F2634FCF00EC8403781025ED6890C4849742706BD43EDE;
precomp_x[68] = 256'h1E33F1A746C9C5778133344D9299FCAA20B0938E8ACFF2544BB40284B8C5FB94;
precomp_x[69] = 256'h85B7C1DCB3CEC1B7EE7F30DED79DD20A0ED1F4CC18CBCFCFA410361FD8F08F31;
precomp_x[70] = 256'h29DF9FBD8D9E46509275F4B125D6D45D7FBE9A3B878A7AF872A2800661AC5F51;
precomp_x[71] = 256'hA0B1CAE06B0A847A3FEA6E671AAF8ADFDFE58CA2F768105C8082B2E449FCE252;
precomp_x[72] = 256'h04E8CEAFB9B3E9A136DC7FF67E840295B499DFB3B2133E4BA113F2E4C0E121E5;
precomp_x[73] = 256'hD24A44E047E19B6F5AFB81C7CA2F69080A5076689A010919F42725C2B789A33B;
precomp_x[74] = 256'hEA01606A7A6C9CDD249FDFCFACB99584001EDD28ABBAB77B5104E98E8E3B35D4;
precomp_x[75] = 256'hAF8ADDBF2B661C8A6C6328655EB96651252007D8C5EA31BE4AD196DE8CE2131F;
precomp_x[76] = 256'h00E3AE1974566CA06CC516D47E0FB165A674A3DABCFCA15E722F0E3450F45889;
precomp_x[77] = 256'h591EE355313D99721CF6993FFED1E3E301993FF3ED258802075EA8CED397E246;
precomp_x[78] = 256'h11396D55FDA54C49F19AA97318D8DA61FA8584E47B084945077CF03255B52984;
precomp_x[79] = 256'h3C5D2A1BA39C5A1790000738C9E0C40B8DCDFD5468754B6405540157E017AA7A;
precomp_x[80] = 256'hCC8704B8A60A0DEFA3A99A7299F2E9C3FBC395AFB04AC078425EF8A1793CC030;
precomp_x[81] = 256'hC533E4F7EA8555AACD9777AC5CAD29B97DD4DEFCCC53EE7EA204119B2889B197;
precomp_x[82] = 256'h0C14F8F2CCB27D6F109F6D08D03CC96A69BA8C34EEC07BBCF566D48E33DA6593;
precomp_x[83] = 256'hA6CBC3046BC6A450BAC24789FA17115A4C9739ED75F8F21CE441F72E0B90E6EF;
precomp_x[84] = 256'h347D6D9A02C48927EBFB86C1359B1CAF130A3C0267D11CE6344B39F99D43CC38;
precomp_x[85] = 256'hDA6545D2181DB8D983F7DCB375EF5866D47C67B1BF31C8CF855EF7437B72656A;
precomp_x[86] = 256'hC40747CC9D012CB1A13B8148309C6DE7EC25D6945D657146B9D5994B8FEB1111;
precomp_x[87] = 256'h4E42C8EC82C99798CCF3A610BE870E78338C7F713348BD34C8203EF4037F3502;
precomp_x[88] = 256'h3775AB7089BC6AF823ABA2E1AF70B236D251CADB0C86743287522A1B3B0DEDEA;
precomp_x[89] = 256'hCEE31CBF7E34EC379D94FB814D3D775AD954595D1314BA8846959E3E82F74E26;
precomp_x[90] = 256'hB4F9EAEA09B6917619F6EA6A4EB5464EFDDB58FD45B1EBEFCDC1A01D08B47986;
precomp_x[91] = 256'hD4263DFC3D2DF923A0179A48966D30CE84E2515AFC3DCCC1B77907792EBCC60E;
precomp_x[92] = 256'h48457524820FA65A4F8D35EB6930857C0032ACC0A4A2DE422233EEDA897612C4;
precomp_x[93] = 256'hDFEEEF1881101F2CB11644F3A2AFDFC2045E19919152923F367A1767C11CCEDA;
precomp_x[94] = 256'h6D7EF6B17543F8373C573F44E1F389835D89BCBC6062CED36C82DF83B8FAE859;
precomp_x[95] = 256'hE75605D59102A5A2684500D3B991F2E3F3C88B93225547035AF25AF66E04541F;
precomp_x[96] = 256'hEB98660F4C4DFAA06A2BE453D5020BC99A0C2E60ABE388457DD43FEFB1ED620C;
precomp_x[97] = 256'h13E87B027D8514D35939F2E6892B19922154596941888336DC3563E3B8DBA942;
precomp_x[98] = 256'hEE163026E9FD6FE017C38F06A5BE6FC125424B371CE2708E7BF4491691E5764A;
precomp_x[99] = 256'hB268F5EF9AD51E4D78DE3A750C2DC89B1E626D43505867999932E5DB33AF3D80;
precomp_x[100] = 256'hFF07F3118A9DF035E9FAD85EB6C7BFE42B02F01CA99CEEA3BF7FFDBA93C4750D;
precomp_x[101] = 256'h8D8B9855C7C052A34146FD20FFB658BEA4B9F69E0D825EBEC16E8C3CE2B526A1;
precomp_x[102] = 256'h52DB0B5384DFBF05BFA9D472D7AE26DFE4B851CECA91B1EBA54263180DA32B63;
precomp_x[103] = 256'hE62F9490D3D51DA6395EFD24E80919CC7D0F29C3F3FA48C6FFF543BECBD43352;
precomp_x[104] = 256'h7F30EA2476B399B4957509C88F77D0191AFA2FF5CB7B14FD6D8E7D65AAAB1193;
precomp_x[105] = 256'h5098FF1E1D9F14FB46A210FADA6C903FEF0FB7B4A1DD1D9AC60A0361800B7A00;
precomp_x[106] = 256'h32B78C7DE9EE512A72895BE6B9CBEFA6E2F3C4CCCE445C96B9F2C81E2778AD58;
precomp_x[107] = 256'hE2CB74FDDC8E9FBCD076EEF2A7C72B0CE37D50F08269DFC074B581550547A4F7;
precomp_x[108] = 256'h8438447566D4D7BEDADC299496AB357426009A35F235CB141BE0D99CD10AE3A8;
precomp_x[109] = 256'h4162D488B89402039B584C6FC6C308870587D9C46F660B878AB65C82C711D67E;
precomp_x[110] = 256'h3FAD3FA84CAF0F34F0F89BFD2DCF54FC175D767AEC3E50684F3BA4A4BF5F683D;
precomp_x[111] = 256'h674F2600A3007A00568C1A7CE05D0816C1FB84BF1370798F1C69532FAEB1A86B;
precomp_x[112] = 256'hD32F4DA54ADE74ABB81B815AD1FB3B263D82D6C692714BCFF87D29BD5EE9F08F;
precomp_x[113] = 256'h30E4E670435385556E593657135845D36FBB6931F72B08CB1ED954F1E3CE3FF6;
precomp_x[114] = 256'hBE2062003C51CC3004682904330E4DEE7F3DCD10B01E580BF1971B04D4CAD297;
precomp_x[115] = 256'h93144423ACE3451ED29E0FB9AC2AF211CB6E84A601DF5993C419859FFF5DF04A;
precomp_x[116] = 256'hB015F8044F5FCBDCF21CA26D6C34FB8197829205C7B7D2A7CB66418C157B112C;
precomp_x[117] = 256'hD5E9E1DA649D97D89E4868117A465A3A4F8A18DE57A140D36B3F2AF341A21B52;
precomp_x[118] = 256'hD3AE41047DD7CA065DBF8ED77B992439983005CD72E16D6F996A5316D36966BB;
precomp_x[119] = 256'h463E2763D885F958FC66CDD22800F0A487197D0A82E377B49F80AF87C897B065;
precomp_x[120] = 256'h7985FDFD127C0567C6F53EC1BB63EC3158E597C40BFE747C83CDDFC910641917;
precomp_x[121] = 256'h74A1AD6B5F76E39DB2DD249410EAC7F99E74C59CB83D2D0ED5FF1543DA7703E9;
precomp_x[122] = 256'h30682A50703375F602D416664BA19B7FC9BAB42C72747463A71D0896B22F6DA3;
precomp_x[123] = 256'h9E2158F0D7C0D5F26C3791EFEFA79597654E7A2B2464F52B1EE6C1347769EF57;
precomp_x[124] = 256'h176E26989A43C9CFEBA4029C202538C28172E566E3C4FCE7322857F3BE327D66;
precomp_x[125] = 256'h75D46EFEA3771E6E68ABB89A13AD747ECF1892393DFC4F1B7004788C50374DA8;
precomp_x[126] = 256'h809A20C67D64900FFB698C4C825F6D5F2310FB0451C869345B7319F645605721;
precomp_x[127] = 256'h1B38903A43F7F114ED4500B4EAC7083FDEFECE1CF29C63528D563446F972C180;
precomp_x[128] = 256'h90A80DB6EB294B9EAB0B4E8DDFA3EFE7263458CE2D07566DF4E6C58868FEEF23;
precomp_x[129] = 256'hC2C80F844B70599812D625460F60340E3E6F36054A14546E6DC25D47376BEA9B;
precomp_x[130] = 256'h9CF606744CF4B5F3FDF989D3F19FB2652D00CFE1D5FCD692A323CE11A28E7553;
precomp_x[131] = 256'h57488FA28742C6B25A493FD6060D936EA6280B0C742005ABCE98F5855AD82208;
precomp_x[132] = 256'hF1133CBE6BE8BBC8DC8DF2B8D75963C2D40ED616C758CDC84EDBC5EB4899447D;
precomp_x[133] = 256'h95083E753301BD787F8989C79065BB813F3D69BFF3E425050F4E04175BBE89C0;
precomp_x[134] = 256'h1A908355CBB756755E576ED29C99AF638668C7B363C8D97362100443BC5C75C6;
precomp_x[135] = 256'hC5922F740BD343D5AA867308FAD97F9F8A2D1F63C5F31DB4F04DF3BEF349B648;
precomp_x[136] = 256'h64E1B1969F9102977691A40431B0B672055DCF31163897D996434420E6C95DC9;
precomp_x[137] = 256'h033B2E76687744ED6C521BAD3333DD37C602F8A7549E9CE7808FB7EA07CE08DE;
precomp_x[138] = 256'h20F18F4C866D8A1CC2A3103317B4AC3189FBF30FF294A75C951473BE45E4F294;
precomp_x[139] = 256'h4D1623C944C9C716A0EB4C685E2A8B9D2DF3465354643BEFD1444176D7B69A8B;
precomp_x[140] = 256'hA901B0DBE8AB292D280D6B36858947854FAAD0A4DD0DA7E2D4AD0FF53DB079E0;
precomp_x[141] = 256'h7E0AF07130218FFD50BD66F4484645B12F42A24F7C80889B3031C9A6EBFC9A70;
precomp_x[142] = 256'h7BA8187E1A7B25A2C185D335440A9038B47F0528546E9DA4EF82AAB05AEBF20D;
precomp_x[143] = 256'h8C050FC34D83B279B6000816E18FCA389767B7960E92677255B84A39D93A6807;
precomp_x[144] = 256'h53B7849A78E4DF8625860583A52499489D7201A2CBF506202A7B8B1BC99C2EC9;
precomp_x[145] = 256'h9BDF9E67A5D0C9956A075A010FE762BEB633500431DEE78EFEBC527E53313B33;
precomp_x[146] = 256'h7CAA72B37A8AB3BD0BAC031A47606F8917D9F42C6EC2D2FB429FD9904A381F34;
precomp_x[147] = 256'h2EF29B9F0982797579C0295FC3F48DB7925D62C75532493DDE16B97E3993D81A;
precomp_x[148] = 256'hDF157CAD95B07875573C1860AE5D02C64029E952EC354E6A9E5C34BE97317FF8;
precomp_x[149] = 256'hDD55C150A29CA526B6182E643B9EB544E651D236B71920E7B15A987016454B1D;
precomp_x[150] = 256'h16886CF46ED42C7919147763063D3256C4D5D39387F0172325B9E4B898227F27;
precomp_x[151] = 256'h6FF180FCDAA3061808E8B306D6F0ACFF27968C22484FF45E56AEAA7B2B60732F;
precomp_x[152] = 256'h03EA4511A00DC2A03EB4F51F40EE677CAA912B5539F685C4F8BCC8EADC395E36;
precomp_x[153] = 256'h0B82CD70DC3DE9EAB38742D8F32DFB8D53E4150A835E54B63C7CCA20F253081D;
precomp_x[154] = 256'hFE2FC3E00074874584EE23BF105A69A606D056F017327D49B7B38B57A196C77F;
precomp_x[155] = 256'h04B90176CDAA369347E8778B12DB9D6EE8B0011446EA35EC845DBF574BB7858B;
precomp_x[156] = 256'h35F382511D34600B4B8C86A9F0DBC9EDDEFC4272F59528A0CD3EC10A5944C6D2;
precomp_x[157] = 256'h1D74B2970311B7FFA1027E26587D3F5BE1D0E9AC3F0111CDF3CC2371722CB94A;
precomp_x[158] = 256'h50A094F309C6F9560B020737B9EC722E4F75D1B7C41593E6F934A68A98450428;
precomp_x[159] = 256'h9B65BB812129157CDFECF12E275EC38C282DBCD914B4810599B0A6D627C63DB7;
precomp_x[160] = 256'h8B4544FC1FDFA06E456C1115A1DC831C85E7F1C5E620ECA51C20802D36A4BC6B;
precomp_x[161] = 256'h6C709880B959EB7C5179B29CC5578FDC6CB2AE13DDCEDE29D5F81D95DE0AB4AA;
precomp_x[162] = 256'h77760B5137BA6A7195D891F794A087A076FC9D67802B81E7085B56773D537806;
precomp_x[163] = 256'h1A8BD7836A0B0C82E9A904A8A8C91A67E23CD4F8EFD625D0DF4C426E7E163102;
precomp_x[164] = 256'hFE217DB659079913FB1E453ED24D91D6A3FB3099E69471D753DB5390864ABC30;
precomp_x[165] = 256'h2504D63754AFD5EBC38F58B65EAD696D07E3ABD748CB6C5F212AED49F5B33B91;
precomp_x[166] = 256'h0B06F702F47B22D789A9BD3F687105C36160ABBF5CC8976B7FBDDCAFDB197B5C;
precomp_x[167] = 256'h803B203BB31F9CF94034EEB931B54480A6F3F99EBD23D0ACBC2128A60D044E23;
precomp_x[168] = 256'h266A9CB4C5F5CEADBB50E5BDA03A7312E52DE1DE8E95A8DCD57289FE0302749A;
precomp_x[169] = 256'hFD8A9D95D80C7AD52599A7AB98163DF364C4C141E9ABEA355D7360BCF84EBA94;
precomp_x[170] = 256'hA7322DF309F28F2359FC339A8B2C80BE6E84ACC5B7B0B8F8F2CB6F26F9DB0A7D;
precomp_x[171] = 256'h82A8C10F336A664963A104DDBF7F0F18BD4C461AEA569FFC82C3C7E4CB052D36;
precomp_x[172] = 256'h9B50D1B68E3BF795007CD12F05A60C266C4EF2B75BA5C516C54784A94F15D6DF;
precomp_x[173] = 256'h3F9083DDC8B423FE7DE3A82281D3056AB8DCB9D7EE82CB806718595FBAE08D32;
precomp_x[174] = 256'hC75C85C1EE17C1A256EFF6BD592666CBC923170659D50BFADBD1074EF2167FAF;
precomp_x[175] = 256'hC5341FEAF8A0F5D3B4D0CF0D2F7AAD7C60EA8E2B3D4B7FB95C68D57698656045;
precomp_x[176] = 256'h83ACDA3E2A8997E0D52BD4C68705DD22220852B7752D67FD8967A03260C2D89B;
precomp_x[177] = 256'h5B8191468B2990745B9C4164E29D594CF1C0D5716C5D39625BD279B30025237B;
precomp_x[178] = 256'h64778122214E38EFF8041796166104E732F5F664D38D77219B89045E2C3B0E6C;
precomp_x[179] = 256'hED4D826AFE5762F4795099099AEE86642B475A9D6DA1017C43D0CB9F1AF12323;
precomp_x[180] = 256'h38B42924419AECC3ACD6F551346FD61A4D82AC2B55F7AFE97A06EB40CD109C4A;
precomp_x[181] = 256'hC3CAD4A8D8BB94A7B434CF70183E8615BB2A8F6224F216E3446AC2E982138911;
precomp_x[182] = 256'h2D408FF4D3D236FD54FAE40DCE3EA9ECD9212E5736591A9E55588E4A54BD6538;
precomp_x[183] = 256'hEE7ADF6D247F25FB76E90CF813F888EBD67423A3A3C6FDAEBAFB7EAA7A33C854;
precomp_x[184] = 256'h2F9457C8A9FFACA13D91151DC4C5E89DDD5D37A37C9A864B7C811F3E01144B34;
precomp_x[185] = 256'hD3F332B8A0F115821CE3478CEFE18DE360120483EF531C277B30C46EB7FEC294;
precomp_x[186] = 256'h183408D338B05AAD3521FCD86EF36DD75F3DDB8666B52F7E9A4CDF1F8E152B91;
precomp_x[187] = 256'h283FEC5DB1145E53BA8F1F0FF9CF89A721FAFFD6C25346863D3956095F40374E;
precomp_x[188] = 256'h0CE7570A4F943CFA413BD249D8E7DBFCEBC73579770FD6DAF54A0DFBDD52FA62;
precomp_x[189] = 256'h7E9C4F19C8F4EC3F1269F648CD919525DF79031574CBEB1537794A4C838FD470;
precomp_x[190] = 256'hE2A9BBE60D5D5BFEA7C7F919DF2309F90BA04F4C722A3EC23BF451B464CB001B;
precomp_x[191] = 256'h504512A43E17EF50E43BF37D42A94990F55E641B1558C265E709900275271012;
precomp_x[192] = 256'h81D1F013A6BB325F4B2D1D51BA72C721859945D8A17B3411CD5CBE87285F850D;
precomp_x[193] = 256'h5B66C2DFC1D2826618A872767E66C33DD90DD51414A3B87CA733383D1D895022;
precomp_x[194] = 256'hAEB5F70E98EC5E38DBD2D544BDBFF8AB99B583D9AF58C597AFAF868820381186;
precomp_x[195] = 256'h0B289EFFE841943B84761E3C67A9C02A557679CA76AD753A707A98212505052E;
precomp_x[196] = 256'hABAE39458B12199E6B0C8360CFD282883F585917E44E1200F81BD356F619291C;
precomp_x[197] = 256'h4A9583A6485B5A5A81AC224A518EB29D1E0F658C8D91B0139419C80955FBACAA;
precomp_x[198] = 256'hD52F630EDBA6F7CB65FCF46544AB0D9EEA236AC1460F17AE3A21010210EBC169;
precomp_x[199] = 256'h0BDC523782C75858F5C50FC052E4C1E9C74A2A6335BCA9BF8D10E1209ADD6A4D;
precomp_x[200] = 256'h44770A338BF0AAB83BB64E476EB6167A88156D168F13CE8626EE0912E59AD087;
precomp_x[201] = 256'hB15E7B322E404AEE319AC20323E366726503108D8EE8E1C83E32D924515E1679;
precomp_x[202] = 256'hA1ED755705225CD0F2C50F758A1C1DF9665AE108D5E0419027BBD9AEDDB00F22;
precomp_x[203] = 256'hE8AAF3616A1BC60FD9BFC43C2C60580F479E9EC9C23A37A23CF8AFB31D918AF5;
precomp_x[204] = 256'h5DC6F8CD2C855E6352A4A4EF6187A6D60759C04338A3DB76C5A3AA37054C20A3;
precomp_x[205] = 256'h6332731167BED8AF68A063EF22AA489CF6563620461AF26A5F1A07CB6B42F3A6;
precomp_x[206] = 256'h8A40D9259A393B382305C2017E8654DBAD66E50AD798A0D3535230F948080263;
precomp_x[207] = 256'hE714710727C7420AF517FD3F9A05B7DEA6A02C8BCC20B17DCDFDEAF82078645A;
precomp_x[208] = 256'h6131291CD95FB87801E42A68553952C29922BCE891C026C0CAE1F69C9661C82D;
precomp_x[209] = 256'h4BC4F845B6764692D0A9BFA81788809EFC5E2AA9DA5003BFB782BCF1D1CA4951;
precomp_x[210] = 256'h45A880A27BBEE9DF29F9BFF5C985F36452865B5D582A201F698E6ECAA2BE67DF;
precomp_x[211] = 256'h6A826A38317C0C8664D6847A220145D1877E5495B21500D3F21F1A0D4AF4F2A4;
precomp_x[212] = 256'h15356506F255F7E96CC8AA1B09DCE5728BD860DE7C6CC75F613E8A34366A23A9;
precomp_x[213] = 256'hF3BC12AEF53D9F5F6B86517802DAC2ECCACFF3A5CCA6443A2B5E1CA0F2B89B91;
precomp_x[214] = 256'h7E3C8C6DFA04A536F7A26EF18B38764922320BEF584533736F728297335C0FD4;
precomp_x[215] = 256'h198CBFCFA0575FC2C161C696D85155FE6943AB9BD6E17223D8844608AD0369D8;
precomp_x[216] = 256'h1E056E89B68CF35A22183C089089B90D5A147CAA780B1FD63AEB1350AFB0E5E8;
precomp_x[217] = 256'hDC7FF9748D827E7EA6173B2F1A646D47D8108144CE7F98FB3FAC729E72FAAA21;
precomp_x[218] = 256'h71B95EFCC4981E0705354BC11CDFBC4836B2EFF0BF8F8EC29A99DA1B2FD28E79;
precomp_x[219] = 256'h43854CAF29DC2BD6C9F3E8FFA25BBA83F6B96121897044AE6876883ADE542B3A;
precomp_x[220] = 256'h02ADFE17090E9F9C708C9B730D5FD084B6EFF990FB87796145C2ECF2D427B222;
precomp_x[221] = 256'hA123452C2B7EAF3115B3A5343B3FF31A09F70C54AE33C620471E3E8227A9D6F9;
precomp_x[222] = 256'h9B89A3C2CA995A8186C1521761348737AAB166AE7DECCA603D06E32CCEC0A6AB;
precomp_x[223] = 256'h64DD7457E7D9D73908E2B9A0DC45272B384B04339ED8B2EDC907964611E9E9B2;
precomp_x[224] = 256'h59227431BE607C6BD327FD714EB71C8720ABBA421C7F550A6B35767D6FA2176C;
precomp_x[225] = 256'h53D765CDADB26E9E1C80DDF199374363843B7D08A7237BDC8C5106EF795FE2C2;
precomp_x[226] = 256'hE507DE9EC16B3BF3523A989C0F5FF6C10452EE909B66FFC16D7B519A57BB66AF;
precomp_x[227] = 256'h016F48C60EB84FB281903B8CB9F60B7A65601D76E2A579835569C98339B4A6F2;
precomp_x[228] = 256'h650471AE774265E3270B513233D12D850BB98E382A3B3AF90CAB6339E1446056;
precomp_x[229] = 256'h15DEA416FA34584FCC90E19D69825FAE348D1BA1FD7AC821559AAC2ABC21DDA8;
precomp_x[230] = 256'hB42B24954F1F70ED3DB900878357BA46EE9D6A07B4F7C751DC5CBA07B05B46E2;
precomp_x[231] = 256'h08E9E4F5C6AEAC311DAB1125DEC9B4606AB10B7E8E250960A17FC57FC0230F83;
precomp_x[232] = 256'h87BE732373BD4B738627FB63BD4D50BFD6F2BB81F804B52829549FE93FE1AC2E;
precomp_x[233] = 256'h43601D61C836387485E9514AB5C8924DD2CFD466AF34AC95002727E1659D60F7;
precomp_x[234] = 256'h341B1580F83071C5365F0BCBBA66AF966902E3942A2560ACA0DAAFA32AB49D0D;
precomp_x[235] = 256'h175E7CB3CE4A3A437C7181E2C79FB15433AC1AA8E56492EB57627171F14DAD95;
precomp_x[236] = 256'h5AD430CC64E61C61E3B3C8482CA3ECAC89C1E4954C80BA98249E45C1307165AD;
precomp_x[237] = 256'h41DCE0D96DACE318988602DF07FA84C1080F0CE3DD7D09F28AEFEFA60DB8B837;
precomp_x[238] = 256'hA5EF449887104DDA103C1DC2520676439AED2D5E0432FE5BA23CC14239961BCC;
precomp_x[239] = 256'h4DA26ECE9AD4600338BDF68B852A2CBE18225F2E2D6D5E626DB57235FB3A9D45;
precomp_x[240] = 256'h6E621E6F53D2408E488D8EB16A19A4F7E9D9558511E6911129DEDC69F98F4763;
precomp_x[241] = 256'hEBAF57645BED74699B57EA758A395A9066BAE20A8F082AB6DA4554D5278BE83B;
precomp_x[242] = 256'hC0F88A71711B632D24B55DBF052B15D2FAA38CA11438C17A6A6FF6353310182F;
precomp_x[243] = 256'h5D9B6C1884B79498C6244FBF262922C6DC1CDDB73CF70AE01B5287B05B5C6350;
precomp_x[244] = 256'hD1D1360F37ED6E69D4F214C6323A53B7E57D759555904016654C49F04E02E21C;
precomp_x[245] = 256'hEFC987CBF1023AF558ACFA1897B1B2B2ACE29A8365674703E4969CCBEE411731;
precomp_x[246] = 256'hF3026B97163DF3BD61B88B7873864480968D1D7B83EF6B0131090FAA18284FF0;
precomp_x[247] = 256'h5D34FF5F123B5B6992AC92C68C9CFF460DEEECF968FF830B5622090D682C5873;
precomp_x[248] = 256'hCBF9BA1794A95247C39DA06584308CC8E0EE591D31A9B0BBDAC67280468447F4;
precomp_x[249] = 256'h920975BA09E2261BBF5982A6B57A73448E7747B8368D7A5379ACACD4C7DCD31F;
precomp_x[250] = 256'h815B2AE46FDCB55D926CDCE82B4F25D0391323123BC180FF33FCF13207EECA64;
precomp_x[251] = 256'h1BB9A6C28E28D4BA30EA86397A4D387E27CA8025DA2319260DE3C454F7E0B16E;
precomp_x[252] = 256'h6F0153FEDFFD83EAB099D29DDDE278F19C05A4BA78EB4C3D34D337C6DA68BC22;
precomp_x[253] = 256'h3454F73B3BEE77A40D00D38471BF555AED23E5E6C6DAE8552E9CB7A91B20258A;
precomp_x[254] = 256'h367807C9A3606B4E1B8C2616AD5280301DFCF68640EDDF02FC59317C230E9A86;
precomp_x[255] = 256'h8EC4FDC39891F6AF1374E06F0C44B81501B8254175FC4909ACBA5941201AF62B;

