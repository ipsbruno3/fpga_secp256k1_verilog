
//-----------------------------------------------------------------------------
// secp256k1_point_mul_wnaf.v
// Scalar point multiplication using windowed NAF (wNAF) algorithm
// Window size: 8 bits (digits in range [-127, 127])
//
// Algorithm:
// 1. Convert scalar k to wNAF representation
// 2. Precompute table: P, 3P, 5P, ..., 255P (128 points for w=8)
// 3. Scan wNAF from MSB to LSB:
//    - Double the accumulator
//    - If digit != 0: add/subtract precomputed point
// 4. Convert result to affine coordinates
//-----------------------------------------------------------------------------

module secp256k1_point_mul_wnaf #(
    parameter integer W = 11 // Change precomp_x precomp_y  with code Folder and change here to fix constants if you change wnaf size 
) (
    input  wire         clk,
    input  wire         rst_n,
    input  wire         start,
    input  wire [255:0] k,           // Scalar
    input  wire [255:0] px,          // (não usado quando use_g=1)
    input  wire [255:0] py,          // (não usado quando use_g=1)
    input  wire         use_g,       // 1 = usa G (tabela fixa)
    output reg  [255:0] qx,
    output reg  [255:0] qy,
    output reg          done,
    output reg          point_at_inf
);

    // -----------------------------
    // Constantes secp256k1
    // -----------------------------
    localparam [255:0] SECP256K1_P = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFC2F;
    localparam [255:0] GX = 256'h79BE667EF9DCBBAC55A06295CE870B07029BFCDB2DCE28D959F2815B16F81798;
    localparam [255:0] GY = 256'h483ADA7726A3C4655DA4FBFC0E1108A8FD17B448A68554199C47D08FFB10D4B8;

    // wNAF "padrão": precisa só dos múltiplos ímpares
    // {1P, 3P, 5P, ..., (2^(W-1)-1)P} => count = 2^(W-2)
    localparam integer NUM_POINTS = (W <= 2) ? 1 : (1 << (W-2));
    localparam integer ADDRW      = (NUM_POINTS <= 2) ? 1 : $clog2(NUM_POINTS);

    reg [255:0] precomp_x [0:NUM_POINTS-1];
    reg [255:0] precomp_y [0:NUM_POINTS-1];

    // Limite de segurança (512 pontos => W=11)
    initial begin : W_CHECK
        if (W < 4 || W > 11) begin
            $fatal(1, "W fora do esperado. Use 2..11 (W=11 => 512 pontos). W=%0d", W);
        end
    end



    // ROM read (1 ciclo)
    reg  [ADDRW-1:0] rom_addr;
    reg  [255:0]     rom_x_q, rom_y_q;
    reg              rom_neg;      // 1 => usa (p - y)
    reg              rom_wait;     // bolha 1 ciclo
    reg              rom_use_add;  // 0 => init_accum, 1 => add_point

    always @(posedge clk) begin
        rom_x_q <= precomp_x[rom_addr];
        rom_y_q <= precomp_y[rom_addr];
    end

    // Inicializa ROM omente W=7 com 32 entradas: 1G,3G,...,63G)
    integer ii;
    initial begin : INIT_ROM
                precomp_x[0] = 256'h79BE667EF9DCBBAC55A06295CE870B07029BFCDB2DCE28D959F2815B16F81798;
        precomp_x[1] = 256'hF9308A019258C31049344F85F89D5229B531C845836F99B08601F113BCE036F9;
        precomp_x[2] = 256'h2F8BDE4D1A07209355B4A7250A5C5128E88B84BDDC619AB7CBA8D569B240EFE4;
        precomp_x[3] = 256'h5CBDF0646E5DB4EAA398F365F2EA7A0E3D419B7E0330E39CE92BDDEDCAC4F9BC;
        precomp_x[4] = 256'hACD484E2F0C7F65309AD178A9F559ABDE09796974C57E714C35F110DFC27CCBE;
        precomp_x[5] = 256'h774AE7F858A9411E5EF4246B70C65AAC5649980BE5C17891BBEC17895DA008CB;
        precomp_x[6] = 256'hF28773C2D975288BC7D1D205C3748651B075FBC6610E58CDDEEDDF8F19405AA8;
        precomp_x[7] = 256'hD7924D4F7D43EA965A465AE3095FF41131E5946F3C85F79E44ADBCF8E27E080E;
        precomp_x[8] = 256'hDEFDEA4CDB677750A420FEE807EACF21EB9898AE79B9768766E4FAA04A2D4A34;
        precomp_x[9] = 256'h2B4EA0A797A443D293EF5CFF444F4979F06ACFEBD7E86D277475656138385B6C;
        precomp_x[10] = 256'h352BBF4A4CDD12564F93FA332CE333301D9AD40271F8107181340AEF25BE59D5;
        precomp_x[11] = 256'h2FA2104D6B38D11B0230010559879124E42AB8DFEFF5FF29DC9CDADD4ECACC3F;
        precomp_x[12] = 256'h9248279B09B4D68DAB21A9B066EDDA83263C3D84E09572E269CA0CD7F5453714;
        precomp_x[13] = 256'hDAED4F2BE3A8BF278E70132FB0BEB7522F570E144BF615C07E996D443DEE8729;
        precomp_x[14] = 256'hC44D12C7065D812E8ACF28D7CBB19F9011ECD9E9FDF281B0E6A3B5E87D22E7DB;
        precomp_x[15] = 256'h6A245BF6DC698504C89A20CFDED60853152B695336C28063B61C65CBD269E6B4;
        precomp_x[16] = 256'h1697FFA6FD9DE627C077E3D2FE541084CE13300B0BEC1146F95AE57F0D0BD6A5;
        precomp_x[17] = 256'h605BDB019981718B986D0F07E834CB0D9DEB8360FFB7F61DF982345EF27A7479;
        precomp_x[18] = 256'h62D14DAB4150BF497402FDC45A215E10DCB01C354959B10CFE31C7E9D87FF33D;
        precomp_x[19] = 256'h80C60AD0040F27DADE5B4B06C408E56B2C50E9F56B9B8B425E555C2F86308B6F;
        precomp_x[20] = 256'h7A9375AD6167AD54AA74C6348CC54D344CC5DC9487D847049D5EABB0FA03C8FB;
        precomp_x[21] = 256'hD528ECD9B696B54C907A9ED045447A79BB408EC39B68DF504BB51F459BC3FFC9;
        precomp_x[22] = 256'h049370A4B5F43412EA25F514E8ECDAD05266115E4A7ECB1387231808F8B45963;
        precomp_x[23] = 256'h77F230936EE88CBBD73DF930D64702EF881D811E0E1498E2F1C13EB1FC345D74;
        precomp_x[24] = 256'hF2DAC991CC4CE4B9EA44887E5C7C0BCE58C80074AB9D4DBAEB28531B7739F530;
        precomp_x[25] = 256'h463B3D9F662621FB1B4BE8FBBE2520125A216CDFC9DAE3DEBCBA4850C690D45B;
        precomp_x[26] = 256'hF16F804244E46E2A09232D4AFF3B59976B98FAC14328A2D1A32496B49998F247;
        precomp_x[27] = 256'hCAF754272DC84563B0352B7A14311AF55D245315ACE27C65369E15F7151D41D1;
        precomp_x[28] = 256'h2600CA4B282CB986F85D0F1709979D8B44A09C07CB86D7C124497BC86F082120;
        precomp_x[29] = 256'h7635CA72D7E8432C338EC53CD12220BC01C48685E24F7DC8C602A7746998E435;
        precomp_x[30] = 256'h754E3239F325570CDBBF4A87DEEE8A66B7F2B33479D468FBC1A50743BF56CC18;
        precomp_x[31] = 256'hE3E6BD1071A1E96AFF57859C82D570F0330800661D1C952F9FE2694691D9B9E8;
        precomp_x[32] = 256'h186B483D056A033826AE73D88F732985C4CCB1F32BA35F4B4CC47FDCF04AA6EB;
        precomp_x[33] = 256'hDF9D70A6B9876CE544C98561F4BE4F725442E6D2B737D9C91A8321724CE0963F;
        precomp_x[34] = 256'h5EDD5CC23C51E87A497CA815D5DCE0F8AB52554F849ED8995DE64C5F34CE7143;
        precomp_x[35] = 256'h290798C2B6476830DA12FE02287E9E777AA3FBA1C355B17A722D362F84614FBA;
        precomp_x[36] = 256'hAF3C423A95D9F5B3054754EFA150AC39CD29552FE360257362DFDECEF4053B45;
        precomp_x[37] = 256'h766DBB24D134E745CCCAA28C99BF274906BB66B26DCF98DF8D2FED50D884249A;
        precomp_x[38] = 256'h59DBF46F8C94759BA21277C33784F41645F7B44F6C596A58CE92E666191ABE3E;
        precomp_x[39] = 256'hF13ADA95103C4537305E691E74E9A4A8DD647E711A95E73CB62DC6018CFD87B8;
        precomp_x[40] = 256'h7754B4FA0E8ACED06D4167A2C59CCA4CDA1869C06EBADFB6488550015A88522C;
        precomp_x[41] = 256'h948DCADF5990E048AA3874D46ABEF9D701858F95DE8041D2A6828C99E2262519;
        precomp_x[42] = 256'h7962414450C76C1689C7B48F8202EC37FB224CF5AC0BFA1570328A8A3D7C77AB;
        precomp_x[43] = 256'h3514087834964B54B15B160644D915485A16977225B8847BB0DD085137EC47CA;
        precomp_x[44] = 256'hD3CC30AD6B483E4BC79CE2C9DD8BC54993E947EB8DF787B442943D3F7B527EAF;
        precomp_x[45] = 256'h1624D84780732860CE1C78FCBFEFE08B2B29823DB913F6493975BA0FF4847610;
        precomp_x[46] = 256'h733CE80DA955A8A26902C95633E62A985192474B5AF207DA6DF7B4FD5FC61CD4;
        precomp_x[47] = 256'h15D9441254945064CF1A1C33BBD3B49F8966C5092171E699EF258DFAB81C045C;
        precomp_x[48] = 256'hA1D0FCF2EC9DE675B612136E5CE70D271C21417C9D2B8AAAAC138599D0717940;
        precomp_x[49] = 256'hE22FBE15C0AF8CCC5780C0735F84DBE9A790BADEE8245C06C7CA37331CB36980;
        precomp_x[50] = 256'h311091DD9860E8E20EE13473C1155F5F69635E394704EAA74009452246CFA9B3;
        precomp_x[51] = 256'h34C1FD04D301BE89B31C0442D3E6AC24883928B45A9340781867D4232EC2DBDF;
        precomp_x[52] = 256'hF219EA5D6B54701C1C14DE5B557EB42A8D13F3ABBCD08AFFCC2A5E6B049B8D63;
        precomp_x[53] = 256'hD7B8740F74A8FBAAB1F683DB8F45DE26543A5490BCA627087236912469A0B448;
        precomp_x[54] = 256'h32D31C222F8F6F0EF86F7C98D3A3335EAD5BCD32ABDD94289FE4D3091AA824BF;
        precomp_x[55] = 256'h7461F371914AB32671045A155D9831EA8793D77CD59592C4340F86CBC18347B5;
        precomp_x[56] = 256'hEE079ADB1DF1860074356A25AA38206A6D716B2C3E67453D287698BAD7B2B2D6;
        precomp_x[57] = 256'h16EC93E447EC83F0467B18302EE620F7E65DE331874C9DC72BFD8616BA9DA6B5;
        precomp_x[58] = 256'hEAA5F980C245F6F038978290AFA70B6BD8855897F98B6AA485B96065D537BD99;
        precomp_x[59] = 256'h078C9407544AC132692EE1910A02439958AE04877151342EA96C4B6B35A49F51;
        precomp_x[60] = 256'h494F4BE219A1A77016DCD838431AEA0001CDC8AE7A6FC688726578D9702857A5;
        precomp_x[61] = 256'hA598A8030DA6D86C6BC7F2F5144EA549D28211EA58FAA70EBF4C1E665C1FE9B5;
        precomp_x[62] = 256'hC41916365ABB2B5D09192F5F2DBEAFEC208F020F12570A184DBADC3E58595997;
        precomp_x[63] = 256'h841D6063A586FA475A724604DA03BC5B92A2E0D2E0A36ACFE4C73A5514742881;
        precomp_x[64] = 256'h5E95BB399A6971D376026947F89BDE2F282B33810928BE4DED112AC4D70E20D5;
        precomp_x[65] = 256'h36E4641A53948FD476C39F8A99FD974E5EC07564B5315D8BF99471BCA0EF2F66;
        precomp_x[66] = 256'h0336581EA7BFBBB290C191A2F507A41CF5643842170E914FAEAB27C2C579F726;
        precomp_x[67] = 256'h8AB89816DADFD6B6A1F2634FCF00EC8403781025ED6890C4849742706BD43EDE;
        precomp_x[68] = 256'h1E33F1A746C9C5778133344D9299FCAA20B0938E8ACFF2544BB40284B8C5FB94;
        precomp_x[69] = 256'h85B7C1DCB3CEC1B7EE7F30DED79DD20A0ED1F4CC18CBCFCFA410361FD8F08F31;
        precomp_x[70] = 256'h29DF9FBD8D9E46509275F4B125D6D45D7FBE9A3B878A7AF872A2800661AC5F51;
        precomp_x[71] = 256'hA0B1CAE06B0A847A3FEA6E671AAF8ADFDFE58CA2F768105C8082B2E449FCE252;
        precomp_x[72] = 256'h04E8CEAFB9B3E9A136DC7FF67E840295B499DFB3B2133E4BA113F2E4C0E121E5;
        precomp_x[73] = 256'hD24A44E047E19B6F5AFB81C7CA2F69080A5076689A010919F42725C2B789A33B;
        precomp_x[74] = 256'hEA01606A7A6C9CDD249FDFCFACB99584001EDD28ABBAB77B5104E98E8E3B35D4;
        precomp_x[75] = 256'hAF8ADDBF2B661C8A6C6328655EB96651252007D8C5EA31BE4AD196DE8CE2131F;
        precomp_x[76] = 256'h00E3AE1974566CA06CC516D47E0FB165A674A3DABCFCA15E722F0E3450F45889;
        precomp_x[77] = 256'h591EE355313D99721CF6993FFED1E3E301993FF3ED258802075EA8CED397E246;
        precomp_x[78] = 256'h11396D55FDA54C49F19AA97318D8DA61FA8584E47B084945077CF03255B52984;
        precomp_x[79] = 256'h3C5D2A1BA39C5A1790000738C9E0C40B8DCDFD5468754B6405540157E017AA7A;
        precomp_x[80] = 256'hCC8704B8A60A0DEFA3A99A7299F2E9C3FBC395AFB04AC078425EF8A1793CC030;
        precomp_x[81] = 256'hC533E4F7EA8555AACD9777AC5CAD29B97DD4DEFCCC53EE7EA204119B2889B197;
        precomp_x[82] = 256'h0C14F8F2CCB27D6F109F6D08D03CC96A69BA8C34EEC07BBCF566D48E33DA6593;
        precomp_x[83] = 256'hA6CBC3046BC6A450BAC24789FA17115A4C9739ED75F8F21CE441F72E0B90E6EF;
        precomp_x[84] = 256'h347D6D9A02C48927EBFB86C1359B1CAF130A3C0267D11CE6344B39F99D43CC38;
        precomp_x[85] = 256'hDA6545D2181DB8D983F7DCB375EF5866D47C67B1BF31C8CF855EF7437B72656A;
        precomp_x[86] = 256'hC40747CC9D012CB1A13B8148309C6DE7EC25D6945D657146B9D5994B8FEB1111;
        precomp_x[87] = 256'h4E42C8EC82C99798CCF3A610BE870E78338C7F713348BD34C8203EF4037F3502;
        precomp_x[88] = 256'h3775AB7089BC6AF823ABA2E1AF70B236D251CADB0C86743287522A1B3B0DEDEA;
        precomp_x[89] = 256'hCEE31CBF7E34EC379D94FB814D3D775AD954595D1314BA8846959E3E82F74E26;
        precomp_x[90] = 256'hB4F9EAEA09B6917619F6EA6A4EB5464EFDDB58FD45B1EBEFCDC1A01D08B47986;
        precomp_x[91] = 256'hD4263DFC3D2DF923A0179A48966D30CE84E2515AFC3DCCC1B77907792EBCC60E;
        precomp_x[92] = 256'h48457524820FA65A4F8D35EB6930857C0032ACC0A4A2DE422233EEDA897612C4;
        precomp_x[93] = 256'hDFEEEF1881101F2CB11644F3A2AFDFC2045E19919152923F367A1767C11CCEDA;
        precomp_x[94] = 256'h6D7EF6B17543F8373C573F44E1F389835D89BCBC6062CED36C82DF83B8FAE859;
        precomp_x[95] = 256'hE75605D59102A5A2684500D3B991F2E3F3C88B93225547035AF25AF66E04541F;
        precomp_x[96] = 256'hEB98660F4C4DFAA06A2BE453D5020BC99A0C2E60ABE388457DD43FEFB1ED620C;
        precomp_x[97] = 256'h13E87B027D8514D35939F2E6892B19922154596941888336DC3563E3B8DBA942;
        precomp_x[98] = 256'hEE163026E9FD6FE017C38F06A5BE6FC125424B371CE2708E7BF4491691E5764A;
        precomp_x[99] = 256'hB268F5EF9AD51E4D78DE3A750C2DC89B1E626D43505867999932E5DB33AF3D80;
        precomp_x[100] = 256'hFF07F3118A9DF035E9FAD85EB6C7BFE42B02F01CA99CEEA3BF7FFDBA93C4750D;
        precomp_x[101] = 256'h8D8B9855C7C052A34146FD20FFB658BEA4B9F69E0D825EBEC16E8C3CE2B526A1;
        precomp_x[102] = 256'h52DB0B5384DFBF05BFA9D472D7AE26DFE4B851CECA91B1EBA54263180DA32B63;
        precomp_x[103] = 256'hE62F9490D3D51DA6395EFD24E80919CC7D0F29C3F3FA48C6FFF543BECBD43352;
        precomp_x[104] = 256'h7F30EA2476B399B4957509C88F77D0191AFA2FF5CB7B14FD6D8E7D65AAAB1193;
        precomp_x[105] = 256'h5098FF1E1D9F14FB46A210FADA6C903FEF0FB7B4A1DD1D9AC60A0361800B7A00;
        precomp_x[106] = 256'h32B78C7DE9EE512A72895BE6B9CBEFA6E2F3C4CCCE445C96B9F2C81E2778AD58;
        precomp_x[107] = 256'hE2CB74FDDC8E9FBCD076EEF2A7C72B0CE37D50F08269DFC074B581550547A4F7;
        precomp_x[108] = 256'h8438447566D4D7BEDADC299496AB357426009A35F235CB141BE0D99CD10AE3A8;
        precomp_x[109] = 256'h4162D488B89402039B584C6FC6C308870587D9C46F660B878AB65C82C711D67E;
        precomp_x[110] = 256'h3FAD3FA84CAF0F34F0F89BFD2DCF54FC175D767AEC3E50684F3BA4A4BF5F683D;
        precomp_x[111] = 256'h674F2600A3007A00568C1A7CE05D0816C1FB84BF1370798F1C69532FAEB1A86B;
        precomp_x[112] = 256'hD32F4DA54ADE74ABB81B815AD1FB3B263D82D6C692714BCFF87D29BD5EE9F08F;
        precomp_x[113] = 256'h30E4E670435385556E593657135845D36FBB6931F72B08CB1ED954F1E3CE3FF6;
        precomp_x[114] = 256'hBE2062003C51CC3004682904330E4DEE7F3DCD10B01E580BF1971B04D4CAD297;
        precomp_x[115] = 256'h93144423ACE3451ED29E0FB9AC2AF211CB6E84A601DF5993C419859FFF5DF04A;
        precomp_x[116] = 256'hB015F8044F5FCBDCF21CA26D6C34FB8197829205C7B7D2A7CB66418C157B112C;
        precomp_x[117] = 256'hD5E9E1DA649D97D89E4868117A465A3A4F8A18DE57A140D36B3F2AF341A21B52;
        precomp_x[118] = 256'hD3AE41047DD7CA065DBF8ED77B992439983005CD72E16D6F996A5316D36966BB;
        precomp_x[119] = 256'h463E2763D885F958FC66CDD22800F0A487197D0A82E377B49F80AF87C897B065;
        precomp_x[120] = 256'h7985FDFD127C0567C6F53EC1BB63EC3158E597C40BFE747C83CDDFC910641917;
        precomp_x[121] = 256'h74A1AD6B5F76E39DB2DD249410EAC7F99E74C59CB83D2D0ED5FF1543DA7703E9;
        precomp_x[122] = 256'h30682A50703375F602D416664BA19B7FC9BAB42C72747463A71D0896B22F6DA3;
        precomp_x[123] = 256'h9E2158F0D7C0D5F26C3791EFEFA79597654E7A2B2464F52B1EE6C1347769EF57;
        precomp_x[124] = 256'h176E26989A43C9CFEBA4029C202538C28172E566E3C4FCE7322857F3BE327D66;
        precomp_x[125] = 256'h75D46EFEA3771E6E68ABB89A13AD747ECF1892393DFC4F1B7004788C50374DA8;
        precomp_x[126] = 256'h809A20C67D64900FFB698C4C825F6D5F2310FB0451C869345B7319F645605721;
        precomp_x[127] = 256'h1B38903A43F7F114ED4500B4EAC7083FDEFECE1CF29C63528D563446F972C180;
        precomp_x[128] = 256'h90A80DB6EB294B9EAB0B4E8DDFA3EFE7263458CE2D07566DF4E6C58868FEEF23;
        precomp_x[129] = 256'hC2C80F844B70599812D625460F60340E3E6F36054A14546E6DC25D47376BEA9B;
        precomp_x[130] = 256'h9CF606744CF4B5F3FDF989D3F19FB2652D00CFE1D5FCD692A323CE11A28E7553;
        precomp_x[131] = 256'h57488FA28742C6B25A493FD6060D936EA6280B0C742005ABCE98F5855AD82208;
        precomp_x[132] = 256'hF1133CBE6BE8BBC8DC8DF2B8D75963C2D40ED616C758CDC84EDBC5EB4899447D;
        precomp_x[133] = 256'h95083E753301BD787F8989C79065BB813F3D69BFF3E425050F4E04175BBE89C0;
        precomp_x[134] = 256'h1A908355CBB756755E576ED29C99AF638668C7B363C8D97362100443BC5C75C6;
        precomp_x[135] = 256'hC5922F740BD343D5AA867308FAD97F9F8A2D1F63C5F31DB4F04DF3BEF349B648;
        precomp_x[136] = 256'h64E1B1969F9102977691A40431B0B672055DCF31163897D996434420E6C95DC9;
        precomp_x[137] = 256'h033B2E76687744ED6C521BAD3333DD37C602F8A7549E9CE7808FB7EA07CE08DE;
        precomp_x[138] = 256'h20F18F4C866D8A1CC2A3103317B4AC3189FBF30FF294A75C951473BE45E4F294;
        precomp_x[139] = 256'h4D1623C944C9C716A0EB4C685E2A8B9D2DF3465354643BEFD1444176D7B69A8B;
        precomp_x[140] = 256'hA901B0DBE8AB292D280D6B36858947854FAAD0A4DD0DA7E2D4AD0FF53DB079E0;
        precomp_x[141] = 256'h7E0AF07130218FFD50BD66F4484645B12F42A24F7C80889B3031C9A6EBFC9A70;
        precomp_x[142] = 256'h7BA8187E1A7B25A2C185D335440A9038B47F0528546E9DA4EF82AAB05AEBF20D;
        precomp_x[143] = 256'h8C050FC34D83B279B6000816E18FCA389767B7960E92677255B84A39D93A6807;
        precomp_x[144] = 256'h53B7849A78E4DF8625860583A52499489D7201A2CBF506202A7B8B1BC99C2EC9;
        precomp_x[145] = 256'h9BDF9E67A5D0C9956A075A010FE762BEB633500431DEE78EFEBC527E53313B33;
        precomp_x[146] = 256'h7CAA72B37A8AB3BD0BAC031A47606F8917D9F42C6EC2D2FB429FD9904A381F34;
        precomp_x[147] = 256'h2EF29B9F0982797579C0295FC3F48DB7925D62C75532493DDE16B97E3993D81A;
        precomp_x[148] = 256'hDF157CAD95B07875573C1860AE5D02C64029E952EC354E6A9E5C34BE97317FF8;
        precomp_x[149] = 256'hDD55C150A29CA526B6182E643B9EB544E651D236B71920E7B15A987016454B1D;
        precomp_x[150] = 256'h16886CF46ED42C7919147763063D3256C4D5D39387F0172325B9E4B898227F27;
        precomp_x[151] = 256'h6FF180FCDAA3061808E8B306D6F0ACFF27968C22484FF45E56AEAA7B2B60732F;
        precomp_x[152] = 256'h03EA4511A00DC2A03EB4F51F40EE677CAA912B5539F685C4F8BCC8EADC395E36;
        precomp_x[153] = 256'h0B82CD70DC3DE9EAB38742D8F32DFB8D53E4150A835E54B63C7CCA20F253081D;
        precomp_x[154] = 256'hFE2FC3E00074874584EE23BF105A69A606D056F017327D49B7B38B57A196C77F;
        precomp_x[155] = 256'h04B90176CDAA369347E8778B12DB9D6EE8B0011446EA35EC845DBF574BB7858B;
        precomp_x[156] = 256'h35F382511D34600B4B8C86A9F0DBC9EDDEFC4272F59528A0CD3EC10A5944C6D2;
        precomp_x[157] = 256'h1D74B2970311B7FFA1027E26587D3F5BE1D0E9AC3F0111CDF3CC2371722CB94A;
        precomp_x[158] = 256'h50A094F309C6F9560B020737B9EC722E4F75D1B7C41593E6F934A68A98450428;
        precomp_x[159] = 256'h9B65BB812129157CDFECF12E275EC38C282DBCD914B4810599B0A6D627C63DB7;
        precomp_x[160] = 256'h8B4544FC1FDFA06E456C1115A1DC831C85E7F1C5E620ECA51C20802D36A4BC6B;
        precomp_x[161] = 256'h6C709880B959EB7C5179B29CC5578FDC6CB2AE13DDCEDE29D5F81D95DE0AB4AA;
        precomp_x[162] = 256'h77760B5137BA6A7195D891F794A087A076FC9D67802B81E7085B56773D537806;
        precomp_x[163] = 256'h1A8BD7836A0B0C82E9A904A8A8C91A67E23CD4F8EFD625D0DF4C426E7E163102;
        precomp_x[164] = 256'hFE217DB659079913FB1E453ED24D91D6A3FB3099E69471D753DB5390864ABC30;
        precomp_x[165] = 256'h2504D63754AFD5EBC38F58B65EAD696D07E3ABD748CB6C5F212AED49F5B33B91;
        precomp_x[166] = 256'h0B06F702F47B22D789A9BD3F687105C36160ABBF5CC8976B7FBDDCAFDB197B5C;
        precomp_x[167] = 256'h803B203BB31F9CF94034EEB931B54480A6F3F99EBD23D0ACBC2128A60D044E23;
        precomp_x[168] = 256'h266A9CB4C5F5CEADBB50E5BDA03A7312E52DE1DE8E95A8DCD57289FE0302749A;
        precomp_x[169] = 256'hFD8A9D95D80C7AD52599A7AB98163DF364C4C141E9ABEA355D7360BCF84EBA94;
        precomp_x[170] = 256'hA7322DF309F28F2359FC339A8B2C80BE6E84ACC5B7B0B8F8F2CB6F26F9DB0A7D;
        precomp_x[171] = 256'h82A8C10F336A664963A104DDBF7F0F18BD4C461AEA569FFC82C3C7E4CB052D36;
        precomp_x[172] = 256'h9B50D1B68E3BF795007CD12F05A60C266C4EF2B75BA5C516C54784A94F15D6DF;
        precomp_x[173] = 256'h3F9083DDC8B423FE7DE3A82281D3056AB8DCB9D7EE82CB806718595FBAE08D32;
        precomp_x[174] = 256'hC75C85C1EE17C1A256EFF6BD592666CBC923170659D50BFADBD1074EF2167FAF;
        precomp_x[175] = 256'hC5341FEAF8A0F5D3B4D0CF0D2F7AAD7C60EA8E2B3D4B7FB95C68D57698656045;
        precomp_x[176] = 256'h83ACDA3E2A8997E0D52BD4C68705DD22220852B7752D67FD8967A03260C2D89B;
        precomp_x[177] = 256'h5B8191468B2990745B9C4164E29D594CF1C0D5716C5D39625BD279B30025237B;
        precomp_x[178] = 256'h64778122214E38EFF8041796166104E732F5F664D38D77219B89045E2C3B0E6C;
        precomp_x[179] = 256'hED4D826AFE5762F4795099099AEE86642B475A9D6DA1017C43D0CB9F1AF12323;
        precomp_x[180] = 256'h38B42924419AECC3ACD6F551346FD61A4D82AC2B55F7AFE97A06EB40CD109C4A;
        precomp_x[181] = 256'hC3CAD4A8D8BB94A7B434CF70183E8615BB2A8F6224F216E3446AC2E982138911;
        precomp_x[182] = 256'h2D408FF4D3D236FD54FAE40DCE3EA9ECD9212E5736591A9E55588E4A54BD6538;
        precomp_x[183] = 256'hEE7ADF6D247F25FB76E90CF813F888EBD67423A3A3C6FDAEBAFB7EAA7A33C854;
        precomp_x[184] = 256'h2F9457C8A9FFACA13D91151DC4C5E89DDD5D37A37C9A864B7C811F3E01144B34;
        precomp_x[185] = 256'hD3F332B8A0F115821CE3478CEFE18DE360120483EF531C277B30C46EB7FEC294;
        precomp_x[186] = 256'h183408D338B05AAD3521FCD86EF36DD75F3DDB8666B52F7E9A4CDF1F8E152B91;
        precomp_x[187] = 256'h283FEC5DB1145E53BA8F1F0FF9CF89A721FAFFD6C25346863D3956095F40374E;
        precomp_x[188] = 256'h0CE7570A4F943CFA413BD249D8E7DBFCEBC73579770FD6DAF54A0DFBDD52FA62;
        precomp_x[189] = 256'h7E9C4F19C8F4EC3F1269F648CD919525DF79031574CBEB1537794A4C838FD470;
        precomp_x[190] = 256'hE2A9BBE60D5D5BFEA7C7F919DF2309F90BA04F4C722A3EC23BF451B464CB001B;
        precomp_x[191] = 256'h504512A43E17EF50E43BF37D42A94990F55E641B1558C265E709900275271012;
        precomp_x[192] = 256'h81D1F013A6BB325F4B2D1D51BA72C721859945D8A17B3411CD5CBE87285F850D;
        precomp_x[193] = 256'h5B66C2DFC1D2826618A872767E66C33DD90DD51414A3B87CA733383D1D895022;
        precomp_x[194] = 256'hAEB5F70E98EC5E38DBD2D544BDBFF8AB99B583D9AF58C597AFAF868820381186;
        precomp_x[195] = 256'h0B289EFFE841943B84761E3C67A9C02A557679CA76AD753A707A98212505052E;
        precomp_x[196] = 256'hABAE39458B12199E6B0C8360CFD282883F585917E44E1200F81BD356F619291C;
        precomp_x[197] = 256'h4A9583A6485B5A5A81AC224A518EB29D1E0F658C8D91B0139419C80955FBACAA;
        precomp_x[198] = 256'hD52F630EDBA6F7CB65FCF46544AB0D9EEA236AC1460F17AE3A21010210EBC169;
        precomp_x[199] = 256'h0BDC523782C75858F5C50FC052E4C1E9C74A2A6335BCA9BF8D10E1209ADD6A4D;
        precomp_x[200] = 256'h44770A338BF0AAB83BB64E476EB6167A88156D168F13CE8626EE0912E59AD087;
        precomp_x[201] = 256'hB15E7B322E404AEE319AC20323E366726503108D8EE8E1C83E32D924515E1679;
        precomp_x[202] = 256'hA1ED755705225CD0F2C50F758A1C1DF9665AE108D5E0419027BBD9AEDDB00F22;
        precomp_x[203] = 256'hE8AAF3616A1BC60FD9BFC43C2C60580F479E9EC9C23A37A23CF8AFB31D918AF5;
        precomp_x[204] = 256'h5DC6F8CD2C855E6352A4A4EF6187A6D60759C04338A3DB76C5A3AA37054C20A3;
        precomp_x[205] = 256'h6332731167BED8AF68A063EF22AA489CF6563620461AF26A5F1A07CB6B42F3A6;
        precomp_x[206] = 256'h8A40D9259A393B382305C2017E8654DBAD66E50AD798A0D3535230F948080263;
        precomp_x[207] = 256'hE714710727C7420AF517FD3F9A05B7DEA6A02C8BCC20B17DCDFDEAF82078645A;
        precomp_x[208] = 256'h6131291CD95FB87801E42A68553952C29922BCE891C026C0CAE1F69C9661C82D;
        precomp_x[209] = 256'h4BC4F845B6764692D0A9BFA81788809EFC5E2AA9DA5003BFB782BCF1D1CA4951;
        precomp_x[210] = 256'h45A880A27BBEE9DF29F9BFF5C985F36452865B5D582A201F698E6ECAA2BE67DF;
        precomp_x[211] = 256'h6A826A38317C0C8664D6847A220145D1877E5495B21500D3F21F1A0D4AF4F2A4;
        precomp_x[212] = 256'h15356506F255F7E96CC8AA1B09DCE5728BD860DE7C6CC75F613E8A34366A23A9;
        precomp_x[213] = 256'hF3BC12AEF53D9F5F6B86517802DAC2ECCACFF3A5CCA6443A2B5E1CA0F2B89B91;
        precomp_x[214] = 256'h7E3C8C6DFA04A536F7A26EF18B38764922320BEF584533736F728297335C0FD4;
        precomp_x[215] = 256'h198CBFCFA0575FC2C161C696D85155FE6943AB9BD6E17223D8844608AD0369D8;
        precomp_x[216] = 256'h1E056E89B68CF35A22183C089089B90D5A147CAA780B1FD63AEB1350AFB0E5E8;
        precomp_x[217] = 256'hDC7FF9748D827E7EA6173B2F1A646D47D8108144CE7F98FB3FAC729E72FAAA21;
        precomp_x[218] = 256'h71B95EFCC4981E0705354BC11CDFBC4836B2EFF0BF8F8EC29A99DA1B2FD28E79;
        precomp_x[219] = 256'h43854CAF29DC2BD6C9F3E8FFA25BBA83F6B96121897044AE6876883ADE542B3A;
        precomp_x[220] = 256'h02ADFE17090E9F9C708C9B730D5FD084B6EFF990FB87796145C2ECF2D427B222;
        precomp_x[221] = 256'hA123452C2B7EAF3115B3A5343B3FF31A09F70C54AE33C620471E3E8227A9D6F9;
        precomp_x[222] = 256'h9B89A3C2CA995A8186C1521761348737AAB166AE7DECCA603D06E32CCEC0A6AB;
        precomp_x[223] = 256'h64DD7457E7D9D73908E2B9A0DC45272B384B04339ED8B2EDC907964611E9E9B2;
        precomp_x[224] = 256'h59227431BE607C6BD327FD714EB71C8720ABBA421C7F550A6B35767D6FA2176C;
        precomp_x[225] = 256'h53D765CDADB26E9E1C80DDF199374363843B7D08A7237BDC8C5106EF795FE2C2;
        precomp_x[226] = 256'hE507DE9EC16B3BF3523A989C0F5FF6C10452EE909B66FFC16D7B519A57BB66AF;
        precomp_x[227] = 256'h016F48C60EB84FB281903B8CB9F60B7A65601D76E2A579835569C98339B4A6F2;
        precomp_x[228] = 256'h650471AE774265E3270B513233D12D850BB98E382A3B3AF90CAB6339E1446056;
        precomp_x[229] = 256'h15DEA416FA34584FCC90E19D69825FAE348D1BA1FD7AC821559AAC2ABC21DDA8;
        precomp_x[230] = 256'hB42B24954F1F70ED3DB900878357BA46EE9D6A07B4F7C751DC5CBA07B05B46E2;
        precomp_x[231] = 256'h08E9E4F5C6AEAC311DAB1125DEC9B4606AB10B7E8E250960A17FC57FC0230F83;
        precomp_x[232] = 256'h87BE732373BD4B738627FB63BD4D50BFD6F2BB81F804B52829549FE93FE1AC2E;
        precomp_x[233] = 256'h43601D61C836387485E9514AB5C8924DD2CFD466AF34AC95002727E1659D60F7;
        precomp_x[234] = 256'h341B1580F83071C5365F0BCBBA66AF966902E3942A2560ACA0DAAFA32AB49D0D;
        precomp_x[235] = 256'h175E7CB3CE4A3A437C7181E2C79FB15433AC1AA8E56492EB57627171F14DAD95;
        precomp_x[236] = 256'h5AD430CC64E61C61E3B3C8482CA3ECAC89C1E4954C80BA98249E45C1307165AD;
        precomp_x[237] = 256'h41DCE0D96DACE318988602DF07FA84C1080F0CE3DD7D09F28AEFEFA60DB8B837;
        precomp_x[238] = 256'hA5EF449887104DDA103C1DC2520676439AED2D5E0432FE5BA23CC14239961BCC;
        precomp_x[239] = 256'h4DA26ECE9AD4600338BDF68B852A2CBE18225F2E2D6D5E626DB57235FB3A9D45;
        precomp_x[240] = 256'h6E621E6F53D2408E488D8EB16A19A4F7E9D9558511E6911129DEDC69F98F4763;
        precomp_x[241] = 256'hEBAF57645BED74699B57EA758A395A9066BAE20A8F082AB6DA4554D5278BE83B;
        precomp_x[242] = 256'hC0F88A71711B632D24B55DBF052B15D2FAA38CA11438C17A6A6FF6353310182F;
        precomp_x[243] = 256'h5D9B6C1884B79498C6244FBF262922C6DC1CDDB73CF70AE01B5287B05B5C6350;
        precomp_x[244] = 256'hD1D1360F37ED6E69D4F214C6323A53B7E57D759555904016654C49F04E02E21C;
        precomp_x[245] = 256'hEFC987CBF1023AF558ACFA1897B1B2B2ACE29A8365674703E4969CCBEE411731;
        precomp_x[246] = 256'hF3026B97163DF3BD61B88B7873864480968D1D7B83EF6B0131090FAA18284FF0;
        precomp_x[247] = 256'h5D34FF5F123B5B6992AC92C68C9CFF460DEEECF968FF830B5622090D682C5873;
        precomp_x[248] = 256'hCBF9BA1794A95247C39DA06584308CC8E0EE591D31A9B0BBDAC67280468447F4;
        precomp_x[249] = 256'h920975BA09E2261BBF5982A6B57A73448E7747B8368D7A5379ACACD4C7DCD31F;
        precomp_x[250] = 256'h815B2AE46FDCB55D926CDCE82B4F25D0391323123BC180FF33FCF13207EECA64;
        precomp_x[251] = 256'h1BB9A6C28E28D4BA30EA86397A4D387E27CA8025DA2319260DE3C454F7E0B16E;
        precomp_x[252] = 256'h6F0153FEDFFD83EAB099D29DDDE278F19C05A4BA78EB4C3D34D337C6DA68BC22;
        precomp_x[253] = 256'h3454F73B3BEE77A40D00D38471BF555AED23E5E6C6DAE8552E9CB7A91B20258A;
        precomp_x[254] = 256'h367807C9A3606B4E1B8C2616AD5280301DFCF68640EDDF02FC59317C230E9A86;
        precomp_x[255] = 256'h8EC4FDC39891F6AF1374E06F0C44B81501B8254175FC4909ACBA5941201AF62B;
        precomp_x[256] = 256'h5CC24A6D4C5B24F914542F91E5FA937FFFA0855151B8B8428729B06A9178A263;
        precomp_x[257] = 256'h83905926C03905C3A9644A6CDA810DD292602A5050C52A219134FC4DE3599E9F;
        precomp_x[258] = 256'h944B097E4721E9DDF8204AC30D3878FAE8FA6C1434AE4822481B29856589B6C7;
        precomp_x[259] = 256'hAB0B4A3FCFB7C134E1CAAF04A63A733117327A1E5FA9030107B5EBBF3423B73D;
        precomp_x[260] = 256'h57A344B5220F2B0EF7BF7FBF05A2E4E71AA2C3D87BF090BCF803DFEE0FE8B85F;
        precomp_x[261] = 256'h6E053E1A800B7C4C51F8C4C95CF0F4FF3608E396EC46188DA1A9263FC8D81AC5;
        precomp_x[262] = 256'h62D764061804717FB30D4A7C7567B54548A289EC7F083F1C59DEAE25CE485CB7;
        precomp_x[263] = 256'hE5DB28F2219FB2AA830CF1080BD2449A5C4D080082D346589E347F31DD29250F;
        precomp_x[264] = 256'h4725B3E9A3D00DE48A53177C9FFF831F733EC89BC2994AB23FE815F109B32729;
        precomp_x[265] = 256'hD0D3AFB6492C72E7394ED9187013E347B036B65EA76E0569BBE9E34641D72B3E;
        precomp_x[266] = 256'h7853E735D717C85797B85654A24ACFF3104143EDCF4B4B4C7869068FC304632C;
        precomp_x[267] = 256'h06DB26B37D4FDC5913A1A01A14C92356EE44E2C97F9D72CA7789DE338EE904A4;
        precomp_x[268] = 256'hB52F0869BB98AF3C0B2F7F5C669FA43E538E400F63A9CCE699AA2EF8EB2848DF;
        precomp_x[269] = 256'h8614DDE11EE6AF03EB34A9E9970FA7C3234152C01384F7E4C1E1F93A0197B448;
        precomp_x[270] = 256'h982A37AE625F6E5B78E71C180F20BDD08B3308EB59D0CAB2DBC20937938C1CFA;
        precomp_x[271] = 256'h6BEA930526B4829CEC99742FC9231C00627A09AF22CA9D9B4081A2FD4C3E703A;
        precomp_x[272] = 256'hB57247818694487E7CC188B336D116B054016A99207319200BA7BD2996583EDB;
        precomp_x[273] = 256'hDE1ADE627BA00E91786F4F5318AC53924DF5A534704EDBB62E0E9E2D997C5412;
        precomp_x[274] = 256'h3738A57CB1721C419F9E465DFB80E1D733720398BC01166DD476D36F3398C0A0;
        precomp_x[275] = 256'h4CAE21C16B2A1239A85575F12DDF6DAA1955FEB8B7502E376940006E7A81885D;
        precomp_x[276] = 256'h4C511A1FBA8A0BE36E37CF5585BCC3A797BFA7EE1BAA60395732FAF8DCC2BD7B;
        precomp_x[277] = 256'hD811D8C4323B43702607C25ADE936C0AC2E4A44B2BA51F8320C5179E745A7E29;
        precomp_x[278] = 256'h101EB5D3B5E5AAFFE39BBAFDF13B5FFA33DB68AE1FB09B0B1CAE25E616C43EEE;
        precomp_x[279] = 256'h89EB1152B8DDE45FE141F21F062FEAD1ECDC7F70EFF8F968DE21CF8B72480519;
        precomp_x[280] = 256'h53D633F3F48EA44D273D8F1E455019A949D95EEB68DE70CDBD1E964D9AD0DC16;
        precomp_x[281] = 256'hDE1069104989110659A94D26B9CEDB646CE3DB4B8398AD1A92F8F95FD8D9BE6A;
        precomp_x[282] = 256'h40ED1E6F0B9EE245AC189A9A7809DA10CC6DAA7B41A163CAF761773C6AF5BEA2;
        precomp_x[283] = 256'h55FAAAEE59A20B9A3784D1719EA529CC1B7AB3A329F26DFAA3B11BD667BA15C1;
        precomp_x[284] = 256'hB51DE64E21CF88AF2180CA1724956D10A95AC607F034FCCBA53BD02BFA8AF3FB;
        precomp_x[285] = 256'h5156B0DCBCD91E824BB235BE9367CF407B8927E8CD874171556F997B7B07B143;
        precomp_x[286] = 256'h3BF51D72060B4973161FAC5588E441A7F1993C06791B6BCD00E11D8E096DD63D;
        precomp_x[287] = 256'hD2971091200881021154F4D3BA6F2DA122FA74C64FAAE05AD76DB7B09AD61FE5;
        precomp_x[288] = 256'hC2EE47CA8E17112FA255A52021FFD30B6D7A3B7E2341526C559B60A9C768013D;
        precomp_x[289] = 256'h559998D69DDCCE0D9E0DA39E96CC4C00C5EF444B561DBAAAE475ADBD3E70B6CF;
        precomp_x[290] = 256'h4B4B02C3E4C8BADDE45305C39721A98D7C1955DD90DCB2F9E9D549016BBAF363;
        precomp_x[291] = 256'hFBAFE7FD7836B42751CF897C5D42897C7650ADE8EE1ED01FE0D7DD2CAAC549C5;
        precomp_x[292] = 256'hCCD306F90C65B8A07884E620B73AC4E681B21BD02A4B219F954DE1B67076C06C;
        precomp_x[293] = 256'hBAFBD838995A691D3B5A870A7847452D9124155DD89A9980820B8D5618195A3B;
        precomp_x[294] = 256'hD125CC3A8073156E0A166AF8FF940A64713D8F37B86919FB157CC380224F458F;
        precomp_x[295] = 256'h7D491F281B5DDABAEF2C6433BE22E42DF2D1BBFD8A7E88668CBF278ECB8187C2;
        precomp_x[296] = 256'h31CCDA339F29123A86C2995C6A9F49796D70A5955079B9616015F07BCDF8C39E;
        precomp_x[297] = 256'h079E64C7F45F91896C92073E71B76FB1E5EC912F0DE11BA7D7439F4A297807BA;
        precomp_x[298] = 256'hD6232EDFFCCB386871EF057B60BDA43F69F422D2DEBCE06C78A31F6A8C42274E;
        precomp_x[299] = 256'h21C0F298B2D6E3A53738FC00C8289458722D78D248A33EA6A7EBB667446E368E;
        precomp_x[300] = 256'h1D1A3D010DCBF799D551621C54F74720EAA2311C3FD9B1D0F4F2CAEE4C3196C8;
        precomp_x[301] = 256'h574886808FA99EDE00CA97D18582A15162E26D5C7753A5614F4BB1DC28E76735;
        precomp_x[302] = 256'hB6DD34D34CE1DFFA4E1E820C4C8BDE9F607194D31C1CE07C9F6FADC89791715A;
        precomp_x[303] = 256'h90F9DED569088772CA2BC8871522DF9B5821DF6C9E20B1600F3504BD4A91D0DE;
        precomp_x[304] = 256'hC55F34E858D193539106E4A0C3002873DB07B2399B10299D260ACC656B2CFA59;
        precomp_x[305] = 256'h6AE44192D38981C59B3F8452C4A2B627F39C16D2B6F525750C5F172256B8ECAD;
        precomp_x[306] = 256'h33A7D639423E1B366A93AD99EAB6444CBD0C251F6CD8B79AE0344EEF6FDCFFBC;
        precomp_x[307] = 256'h48471331EAC4867028FA6642A76CA6C53380C1D90F52A4B2EA640D47F159AF0A;
        precomp_x[308] = 256'h0565AC399AE731C04CFFAAB743D24B7172DEFD79BEB8CE86D46012A5C2587917;
        precomp_x[309] = 256'h964838B53B6C2B7D6A8D017D0C5A32FC995490946DCBF773EAA7085C98314C0B;
        precomp_x[310] = 256'hBC00DA907B8D078B9D83522DAE548B146F9BFF0D02EF887C4AAE2F1EC4EB88D5;
        precomp_x[311] = 256'h1A59F85500F89F0CF13DD8AE9F5E550CA2082BB327FB111D075455ABDBA7BEA4;
        precomp_x[312] = 256'h7A3B611BD3BFFC6AD450816245695024452706A3279A6FDAD88598A54ECCC764;
        precomp_x[313] = 256'h2FED55779CBE0A5A786FA95B5C56E27AA0A1CC2851112BEF4CD5E1B7015D6D91;
        precomp_x[314] = 256'h267AD217952EDF65673EFAEA6BEBB44B018326DDF1B36D02F0154A0D774A9558;
        precomp_x[315] = 256'hEB6ED62C239B99C86978CCECA5F321450E0D341BCA7EAB106FA05EE17F6687E8;
        precomp_x[316] = 256'hCA5CF17CE03D214F0B4EF33C41686C4F5087A59BF88CA7B10891094D430A9E5B;
        precomp_x[317] = 256'h4C7BC29CACF0642E63F035ECA93E6B6CC82F21CF46623A2FE4C7215E51E82F7C;
        precomp_x[318] = 256'h57CAB8E9B42289F0503E50130ACF4DD7797831842389FD2080B61BC3671058E3;
        precomp_x[319] = 256'h3C2BF23DF1120C34DE813A82A56843F5ABF3D272ED2E6C2753FF63109BC4823E;
        precomp_x[320] = 256'hC010A9AC83E0742A0D3348DC3DCFDDD234170AA228D36856D8581B1A0EAB38D2;
        precomp_x[321] = 256'hA4ABD9EE548BA4680E4CB632B3D9C8A94F1B773FBA3A96605504593A92071994;
        precomp_x[322] = 256'hDC02C852EFC115F1C5C08540DECEFFE5D68B82E599B787115A7A333DE8DDA172;
        precomp_x[323] = 256'hEE4769E8223822FFC28A5A4B5F29FD7C0A54FC8172175CAC1B6DB5A291EC57C8;
        precomp_x[324] = 256'hF3006C1D34910C0FD435A6DECF088C382CF990CF3124F2ABB11D2727D93EF066;
        precomp_x[325] = 256'h7CFB203D07BF5669129F0A3E325C3FD6B1B9C8044932F0F3794B93571E7313B7;
        precomp_x[326] = 256'h0CCA3CE036E0099309D30BE8E70455ADEFEABE7183AEB206A324D0EB32312C0A;
        precomp_x[327] = 256'h9FB6414881CD5C2782DA071C01F98D71D9815FD22389D212C66ACE660AB0D9C8;
        precomp_x[328] = 256'h01DBBEBF03E3D45910D39DE232560B4DEB5D2AD806AA1542C2C070B651558B25;
        precomp_x[329] = 256'h7751D21992F474217742856B04C84D415A890EE924185E215A210A3FA46BB5F7;
        precomp_x[330] = 256'h39A849A05B189C3E20782983ECF664B1E7B89C964E11D73770797FCAECF36A2D;
        precomp_x[331] = 256'h67E56125B29CED20F9F95522D412D67C80E3D628B8BFDDEA768117CBE79B25BB;
        precomp_x[332] = 256'h0A51AEDA02F7D59DD31EEC20E95839F6ECDD01EF529327BB5CB229B7B78F1525;
        precomp_x[333] = 256'hC980693E73A1CB46F5EB71B773B00389F8BCB36FFB489E7AAAE64C236AC1745D;
        precomp_x[334] = 256'hC78DF930BCF54C1C28E27AAB2975E9F394167BD2948D47136B17A3740A1391A9;
        precomp_x[335] = 256'h9A75F7BCC6D2F3A9E6168EBC8F7F1E50A998B1E4E67316E5FB242FC46D284089;
        precomp_x[336] = 256'h76B2131ADB0BB3E7DB48277D95CE73E47EBA1E7CB6F801C0D20B71A38B6E6224;
        precomp_x[337] = 256'h218983614EC5971DF55F96C93DA89483CDCC4C46DEB8DE68F32A42B35C1384E1;
        precomp_x[338] = 256'hAC0B0A494E9D180D101DBE1CA528FECBA08449A6CF5D82A9AA14F875E3DB8ADC;
        precomp_x[339] = 256'hF869B58C0851A65FBD6D332975F596A29D1A78CDBBF04A1B6DCA6C2730E04625;
        precomp_x[340] = 256'hF74F02DB2406250F8984A5F2273C63EDA640A43A8E7D72AAECF78D6EB9544C3A;
        precomp_x[341] = 256'hC0613EB61D6755EB2EBC9284A0AA69D288C390504B7E869FF3D943AA067EA65D;
        precomp_x[342] = 256'hEB66FF9860BA08A63C0FD8C47117AEB0AE0DBF63524307A7EB739F08F31285DB;
        precomp_x[343] = 256'h3A7108E6A1256061FC25D58BCA534602E41C6B15156C15B871A516F0EC4A861D;
        precomp_x[344] = 256'hD17E3A58C83169D133EE73717B205F2CEA1A2FF34E744958949E9403B8F89D5F;
        precomp_x[345] = 256'hD6E32892CEFBB8ED14350CBF2618E2FE98CAF6D4F7679385FFF36BAB0BF6541C;
        precomp_x[346] = 256'h318D49FF60E900AE6E8E2182F38EC00682DDC8AE93AA629186D5DDF80AFFEF75;
        precomp_x[347] = 256'hFD6F9E301772DB8BA68EA5AEB585ABBDC075E72B68D6F67C5A2F814498CF6346;
        precomp_x[348] = 256'h8FE25B38A2C74761A90ED08D4BCE768CF074282AE9560D31566AE43A182DDD36;
        precomp_x[349] = 256'h37CF0ED288ED8FEF4AE17BCFF6BFB8153E12BAB2A46D7E5D2E6FEB999793BEF8;
        precomp_x[350] = 256'h688C206106B9D0C876DEB812B60000E8ECA0E04F531ED1E00915844207BF403C;
        precomp_x[351] = 256'h4B4CAAAAF5399535D822371D63965216D1B53584D89A84E9D868395A70B3D804;
        precomp_x[352] = 256'h6F5ACBC44135DA60758ED9A518B39B5F47CCA39824E20E561444DD52E2FA1D2E;
        precomp_x[353] = 256'h79D2D4493DFFCB916FDA527BF8B6B622661D6F23738288C6CE94313DC267FC42;
        precomp_x[354] = 256'h33A8E87E246B7B9C9C77A6B07CC67D41F3915DBC02180118C0800B33F9F95524;
        precomp_x[355] = 256'h9A169132F3887DF820561A7AE4BD54613235DDB20FBA7A193F4DAABA79868E95;
        precomp_x[356] = 256'h790B74F48405CE3F9ABDC7E90439F2F5C859989E2CA5E6FC290461048783AC42;
        precomp_x[357] = 256'hE2A3D0CFAE1FC2D987CAAEB69F32FCD695471785F524E438B5487AA372F9E49C;
        precomp_x[358] = 256'h0CB30C435992C19576D372B196F2AE68CFD2653E63E3BA7A2B3C21EC960BCBEA;
        precomp_x[359] = 256'h1FAEDC95D6310BEE6298FFB16FB3E6A3296CA66B7C995D2DFE92438110E8B46A;
        precomp_x[360] = 256'hA646CF5A2BE8C1D13F05410CED51B3F58E93EA531E28BF318F6C750B52B3E8F9;
        precomp_x[361] = 256'h3273472718537D38E9B8C397A5CC322D1C77C0C615EDED39DCEBC020DEBE2205;
        precomp_x[362] = 256'h16A1A7180855A212C068C095D930A2709906DD22E7DB3F4D4CE2F393D572827E;
        precomp_x[363] = 256'hB4BF4D145DE2557133694B8676166E90EEB1EBF84A7402E9A61AF4CF23687596;
        precomp_x[364] = 256'hD4ED67A9CCF4665E418A0DE08D9380CBFC311413E90A964BBF367B9B0B892630;
        precomp_x[365] = 256'h8AD256F19F413EF20EAE906F0C1C2CA444D5DFDCF916D366B32F1F47F54FE70D;
        precomp_x[366] = 256'h8DD3E2FAFE55B5F1F13723E01A5587B9C67D22EE21F1F62F07F62A1531F17F8E;
        precomp_x[367] = 256'h44FD9E282A8E30AFAC34DB01A7B0E93903C13917554D9A678E577A5D04B3D0F6;
        precomp_x[368] = 256'h5D249A024464ED65831D2AA9C9645F462DB7C9F4E5A46477746B1A7188B7AA42;
        precomp_x[369] = 256'hD98EB4581EDCD51D465E123CD891C481DDD18B540B9408CA85AC47C80E10FB23;
        precomp_x[370] = 256'h2F12C36919A2AEB62132134D2E85150F6EDB486E9D672EB5876804D644DB6082;
        precomp_x[371] = 256'h4D9496847099C9F8421D35DFEBCE57AA713260348F07E3E6F03017C3144B4624;
        precomp_x[372] = 256'hCF1DB9105E95F1C8E360B39A752AB17E0FCA8F24D9DDC8B2A9768700E2AF2466;
        precomp_x[373] = 256'hE71EB4257D2FFA8AB79D63A242C67585D4B1747F05B27F22A9EE42846AA62B85;
        precomp_x[374] = 256'hBCD987D30B2575F43BC5C3E1B4A299BF21C58B6CA27EBB218F9882AB30559887;
        precomp_x[375] = 256'hB74D5CF748AF7162395D2D5E8A69F7407A2BEBBA69564042EA9C7E34B1F8CAB0;
        precomp_x[376] = 256'h46F3DEF59835C9AE1A7B3B13A920BEA9E9BC12EE633B3EDC57251B723560837D;
        precomp_x[377] = 256'h8D3418FDEB3F0968DE51F4D7CBB60299A50CEBA41915D8B65774CFB77667D572;
        precomp_x[378] = 256'h98CB0F094510695D78A0A672EB67253A30F4327B7864FBCF529CF212AD6F7C10;
        precomp_x[379] = 256'h96045E4C0CA075FC4A5383F3F03DE105A34C7C4CB030CEFFB58B98E12B39A3CF;
        precomp_x[380] = 256'hF262E89142ADDEF8CBA26A9CAD779761C3F4B3E55990A93E703BF56A99CC6030;
        precomp_x[381] = 256'h0CD79C02EE1753365F9F7900BE51BB2BAD75EF813C6C56347CC717DB156D17FE;
        precomp_x[382] = 256'h28B4BF225B1D40DDE0122E03E630830AD9BA4629CC51C9D280A225F948F858F4;
        precomp_x[383] = 256'hF018F2067DD55DF39C53344BC6128A5FCC765C36C7B0BEA016C8465CC6ED2FF7;
        precomp_x[384] = 256'h496968CF08086D029A5DD5C74F47CBDA7F661EF1488B394218ED886C424A7A13;
        precomp_x[385] = 256'h242D4C59E9113B7768E4857493600DA7B984355CA1D079498921016B22EFEDAB;
        precomp_x[386] = 256'hB6B804CC1A1A59D384C4AFACC5E5050F466280BCD5AB15861D20F4DD1385E8C7;
        precomp_x[387] = 256'hDC30A3D07ECC5FDD38B8048AF281024B46904B2D2A4C51CA0D1B49B71D918A4E;
        precomp_x[388] = 256'hE1FE434D345BF33083ABB6280F4F44AC5FB22934977813C20C015F2B43D3FAB8;
        precomp_x[389] = 256'hA8ED88DAE08AC5E2AFBE4A40EE77564582C2F513CFD72060BD1FD5D176FB8D08;
        precomp_x[390] = 256'hB52CF828DE1E9CD7C95C083EEC50D2288E770713A0E2543F76FA57902C7C6481;
        precomp_x[391] = 256'h702079AEF76D9BFDCCB957A94AAD93FCB1297C54D634978E4DC78292161D5E83;
        precomp_x[392] = 256'h4638D4D18E9DE1CEEF4FE8CBDB4378E23ED3DCB9513CC9A0DD73EE2EBE57BBF5;
        precomp_x[393] = 256'hEEB34EB75FACADDED561DC5EE3D0A039D98E4880910439CBECFB22D93B386BFC;
        precomp_x[394] = 256'h07F2C6E5BECF3213C1D07DF0CFBE8E39F70A8C643DF7575E5C56859EC52C45CA;
        precomp_x[395] = 256'h6EC767221EC5D27CF7E11064D4F8B0163CEA090F6A950F818562330323E53647;
        precomp_x[396] = 256'h98F6F69D320D5ECA01F184B0378F67CDB44A707AC5B2AF5499E9F8A4524DEA7E;
        precomp_x[397] = 256'hCF1EF44558B82C765D77AC998C0170C92D3086682D9ED7AF2961CF055B47E390;
        precomp_x[398] = 256'h10E01651EFA26F2EF88CC5C10594F3789AB62B825A0875AA37C280A18C6F07E8;
        precomp_x[399] = 256'hB94E2FE041CE209B6EFD77D7449831300AF90945120B9A5805427966E93EEE4A;
        precomp_x[400] = 256'hCF9E7D02C671A9EA145D233E244D8AF66D71CC34E17F2CCC1225D2B316D41154;
        precomp_x[401] = 256'hDA3A3C2994AD3B91319D18EBDCF4B934DF8E4F2BE052F4366D539AFF4BD48BB2;
        precomp_x[402] = 256'hAB8128182B80378BD914C9FCD2831F30A0A095C9D0E52450D4BA27B0F1EEC101;
        precomp_x[403] = 256'hEA5B82A2BF02CAA5D5D64391C0965C53F0EDD967F8DF94AB831408F7E5C4977A;
        precomp_x[404] = 256'h50605C0BAB201D7D03DD618BE3DA2D29318AEAC17DF58D2CA95B8FBCFBE70FA2;
        precomp_x[405] = 256'hF76C50B66D7DCACEF45409D8854F79B651356661108B716831B58B25EA1191DD;
        precomp_x[406] = 256'hDE5053BAD716047CCC2367DB272E4E11413126902BD79B32F6D3D95993260E7D;
        precomp_x[407] = 256'hAD3E719F180E946B1B98A332BDE18E54437F1A240949D7121AFF7C8DFA06499D;
        precomp_x[408] = 256'h270A02345560AF6B6310C867332F8B79839A3AE76E2666ECB46C840CC36BAE4B;
        precomp_x[409] = 256'hEB5ED17E3027C9C4C87FFDB294A84FF725BA2B5B2BF72D30F98334EE68624621;
        precomp_x[410] = 256'hB9C11DF28A0B98CC623F4E8075ACD469FB1F6621A7572D6A7BAC135C2CE0A5DD;
        precomp_x[411] = 256'hEED1704380ABE259FE6611066EDA0408F60F13993C49A21CA8A6310CEBE74B5C;
        precomp_x[412] = 256'h8E4B0F6F5F5B9CF468E5524A4ADF62B68C68E3105EE374C25265000C53AA97A7;
        precomp_x[413] = 256'h77AE21BDFC6596B9AE85CE9C93112B1DA7F393DA1238D76E90CF59C8CAA5EBBE;
        precomp_x[414] = 256'h1D379CA871C02EF459A8BD35F506626592922533F0503999E16D6B07DBD2346F;
        precomp_x[415] = 256'h625017F328FC16AE993671995F02772A5C7EA7217D47C296CBAD670C3FEF1CCC;
        precomp_x[416] = 256'hC7A4FE496BDC35093AE3F508D43877E8D1019D16740A5EB78EAA72B80638412D;
        precomp_x[417] = 256'hCFF9F83CE8F9C4EF3E80102CBC48C409B65C6166B74F052FA5628348B2441D3F;
        precomp_x[418] = 256'h8402771045B8C295C938AE98A9EA11DC2FD23AE57ADE6EF82C60472166700541;
        precomp_x[419] = 256'hF7AB1330E00CB9EC061A346BD8F5522D5E304A4EA94F84AFB5C706140D2E0D2C;
        precomp_x[420] = 256'hA7C84E192303B7788C1A4D5B786C9829D0DA4DDCC13F692C7851884C6FD4E618;
        precomp_x[421] = 256'hB8B0C884A680DAC0363BC55AFA677A72C65F413907F5CDCCF199D80DAC98C43A;
        precomp_x[422] = 256'h816EC443D05761355A3BC33C1DB4A179C5BEF98E943AF8DDAC250482A65E0DF6;
        precomp_x[423] = 256'h8DED2103823D07D533FBA24F7FCCC47CB101960F3B717FD2AF39D49AA91E28A0;
        precomp_x[424] = 256'hB1C4B39CE874D478BFBDF9E3CE8C31650FF4F7C4BEE20C874849AEAAD0D6260B;
        precomp_x[425] = 256'h7D5BCE3BE5953EB3A17F657CFABC8209F011BCF27E10B90D0E75DAD9FAB2C971;
        precomp_x[426] = 256'h2AF5111A422AF2CD14E7717FBC7171C4096AF1788B229497A54D2B874C00F285;
        precomp_x[427] = 256'hB46E29C06DC8DDEFF8BDFB65F4043B61FE010DAEA2D0955DC81A7B49637AF766;
        precomp_x[428] = 256'h105786D3F44EA40F71EB3BD5339CD514AEF6D8FA5923B4A5089B219CFBA6B1EA;
        precomp_x[429] = 256'h1F3C0C81BE856E3018934573892CEB22D2D2D8EFF08B78575C624F4816ADB23F;
        precomp_x[430] = 256'h16DCBAE3A95A95FA0912484FF833BA0EE437876BF16F9C9F5ABF46AA468BD2B3;
        precomp_x[431] = 256'h114BE56CD6723C8F924FF3C0F5EDABC6E42314A649EDBFFF1C794438DAE70726;
        precomp_x[432] = 256'h8D0CB2E601F98472E169DBAC7F5BABFF51766B3A8D74E17D747B7EACD903FDAF;
        precomp_x[433] = 256'h5B420754188C82E4DB72F3A2C804969134E3B43E484B45CAAB4727F531714DB3;
        precomp_x[434] = 256'h91E3761D95761D968D856A72800FE0B59F01C62E1CC446ED18C1B58F88CBF74B;
        precomp_x[435] = 256'h31380B83DC77E5F29C2F55480ABE052A016E0F1F02D8AAD35B05D29C5C1A4655;
        precomp_x[436] = 256'hAE40198CBCD54264904B44C7C90195538F3F3727A0C9639A764CDA80B21EDD27;
        precomp_x[437] = 256'hF4729787ABEAC0F1249B1D3AC19BB0255764A854727B415F73E24C88A8A981C8;
        precomp_x[438] = 256'hF92F02B834148934F7059B617E84D0A6F52D3B8C0A7D7B69CE4C81757ED5884A;
        precomp_x[439] = 256'hA2BED8AAE93BD6820BE8CC4DD1F84FC29EFE4022B2B0DEC49ED3CE177CC93363;
        precomp_x[440] = 256'h5A42CFCD3D1811D199B09DC809308134CF6219E2E029598E899418F9B7AF4724;
        precomp_x[441] = 256'h1D27AB0567E8BF19323F1ECA441750852E768A6BA143678940BA2B945B0E530F;
        precomp_x[442] = 256'h592BF85922C05BF44B42FCF6E4CDF3FDBBBF8088B7263D319BC749146EAB4326;
        precomp_x[443] = 256'h66730A705AE3DAB8BFC01F4ADEEADC410D4DF156D03C4FCF1DD9E16F009359D5;
        precomp_x[444] = 256'h3D002600532420AC09FB246D84E485601CE6897B979491AE07C5914EDBB7FE83;
        precomp_x[445] = 256'h0D42AE362B5DD22FD2089D37D22E2C2A750395AD710AA1C061ED427543A24487;
        precomp_x[446] = 256'h37C761CA486FABFD000B306DC18E9074409E101E5BDD1670EDEF1253AA253743;
        precomp_x[447] = 256'h4E672EF8BBAFBC8EEB819F3715AC0D6C2AFA9781A197345B2889ED0AF3B0E788;
        precomp_x[448] = 256'hC1F2943B23C07929E9C635AE66F6294908E1DF12F35ABA68ED8791D68FD51FEC;
        precomp_x[449] = 256'h3DF2461E739CD98472CF10CDF663E651351E826D7AFDCFFCE17602AEC0370BE6;
        precomp_x[450] = 256'hD4D3D528F98B92D5F4C4ECFBAB60FD8550F123275B63B3FD5518C1F3D62A82B7;
        precomp_x[451] = 256'hECD8399B4AA3368F1A7A411363FF03A7AD6448470E225108B3EE7D021209236B;
        precomp_x[452] = 256'hD5990BE57E6A0DA90333354AFB344D59416D1A70785CDAE38C332E09CDF78722;
        precomp_x[453] = 256'h7598AB651D8CED00AF3D5978661D801EB57E9089287BD74F85EF042A90374B1B;
        precomp_x[454] = 256'hFD071417B12D2D31852048B761C5301BBE088CFD98EBCE7D7E0922CF41F694E7;
        precomp_x[455] = 256'h5A5B4990E290868AD1D571AC8E9347F2B1E513BFCBC2B8D15E56CE012B72CA0E;
        precomp_x[456] = 256'h93DEEC243CD4F14642F5A415F6EA6F3625C900815F3D20F59728C056FDE7F2BD;
        precomp_x[457] = 256'h9224D17BA65AD967969104C93068D4399C9BEC7E7613A602F5C9917E46DF82B6;
        precomp_x[458] = 256'h851ACC9124DDFF9C14CF054B87347A71CFC916376E5591890F0551433B79C38E;
        precomp_x[459] = 256'hFF6C1303B7C111C5087E01EF44829510EFF0A612931F92122B71075F2CEA4D96;
        precomp_x[460] = 256'hF23BD9F055E7BD1D433FB51EC8B6ECB60FD5014F4F4CA9D06A4BC636435FDAC0;
        precomp_x[461] = 256'h9D622C56EA6D5D197B823E601BBD4AF01FE070F9391BB5642A05527A49F46FF7;
        precomp_x[462] = 256'h9494EFE4CFF5D5E76394B67C407B99612915AFDE56933B80370D0ADF2F020C13;
        precomp_x[463] = 256'hA8E4D7BAFFBC52FC00A8CB6C2938A01CE028C25997403268DBE1600A952E1A86;
        precomp_x[464] = 256'h83841F64938E460FEFF191AD4D72D7A5203C01AF1519CDF1F17C3BB5E4927AC5;
        precomp_x[465] = 256'hEE8974D95EF03F8A860DCBA67B597FB2AF2A2DF6950AEACBD623C883020612F6;
        precomp_x[466] = 256'h68E88D8C23616CA3B136E5FA3427628DA92DDE6B2691D857B2D01A60B6579606;
        precomp_x[467] = 256'hFE34DD8AC62EC8B620DBEA7944CCCA40CFE6AB5ACE3B2E7C50AC589A9522345B;
        precomp_x[468] = 256'h423A7A9CC0F81489AAA62479C131736809989366FD18BFF7F6A5F2358251BC1F;
        precomp_x[469] = 256'h7FA60BF97CBF54FFE61BB840B2E08D910FFB0EB4727C0E730ED4F157AD0B98F4;
        precomp_x[470] = 256'h9E53CB0EF1EDDEBC77EDF8A66917F9158294815D0EEF898CF1E7743360153A66;
        precomp_x[471] = 256'hADF93641C616C67799B44AD5354332C01404718E8EC91E9631E695523AD6F119;
        precomp_x[472] = 256'h0701E3EC485DB367B0687DDB2BE15F4B5B6242C4396F6F0C9726ECB6474E4CA8;
        precomp_x[473] = 256'hD8FC5BA5D3ECAA059E9A7E042C52500AD513645E06149E84AAC0D910F8CCFEFC;
        precomp_x[474] = 256'h7BC88F9A8279FFB70658A186FAAA5F0CC900CB9D4A33B8DCC9EEA83EFF71398E;
        precomp_x[475] = 256'h8578D5310BC79E1F6E219BC77F2172A3E5FB92A5EFBF99190F46EA116F5EF0E5;
        precomp_x[476] = 256'h98BC22D73EA2661B545EB5F437E1CC0AD412402044BB90935CDDE758A8020A62;
        precomp_x[477] = 256'h7FCF821E95D2176DD088106CA5BF08559980F265EA3C401AACA44B0AD5E8EE10;
        precomp_x[478] = 256'h898A39B9D440EF05F87E195B6A334F9367ACD67A1FC76CA8316292EA0216A5F1;
        precomp_x[479] = 256'h3EE974A28918C2160A9624801F18BF9A87D6A62783323E3CBF138BF43F2192A4;
        precomp_x[480] = 256'hBDD10D2FDE76DF349AB753EED06C12519766BBF42FB610A57DDC3F364047C14A;
        precomp_x[481] = 256'h2C179437397841244FF9A4A0EB9FF292477A5148C4176B23C000A1CE3BEDD63D;
        precomp_x[482] = 256'h282EF30EF2D61D136F71E6DF6EE97EBDA83036A32D3CD84136289798B3E71580;
        precomp_x[483] = 256'hA42B4D5542ACFA7CB54AB3D50EE0BEBD085BF6EADB138EF71EA38C73899EFF23;
        precomp_x[484] = 256'hB23ACC64C5B00C8F4B580D4749589559A06FCEA575F3D38B1A02251EFF7EF00E;
        precomp_x[485] = 256'h0942DCE696AEB0634681CE7A407516E989DF029CECC77023411A628F75885EA7;
        precomp_x[486] = 256'hB8A6A2B952194EC08238E4DBE71EB94823E64A94E10EA0E1610465AB88392D16;
        precomp_x[487] = 256'hA36D3369A1EE05F7B1FDB083EA614CB6F15FEAC417A416D90CC83FC20868FC20;
        precomp_x[488] = 256'h4EA301083D711AE6FFCCC89B9D6FD4D56F03BD68F4508CC0EBEF5E43088DDA1D;
        precomp_x[489] = 256'h202287161C1C89C764742E62E427B7120FEE118F406A175ECE2F424E2AFFDC55;
        precomp_x[490] = 256'hD3C072FC8E4BF1605790D4296120612395BE9092F166784CF5ADB7E86070D20C;
        precomp_x[491] = 256'h294DAC7CE307FA7CCF0E8F3428A354D294003DBDCA763DAD3E6DF60E0530EC82;
        precomp_x[492] = 256'h3956CA5CC09FE8D9E4042A8D67B276FE225DE609EA24575C7075D9AC4E732FAE;
        precomp_x[493] = 256'h24D2E396DA144B48E736EB06849401754F4109D66D87A9E697EE82BF91FB3DEF;
        precomp_x[494] = 256'h638D4042F16E5C07FCBF9619DD9C2F91188528893E12CD3AB49E2B9B99A2AA5E;
        precomp_x[495] = 256'h0F91AD5BA99972BABB323A1FD3032E1D94202D8863680C5CD7D678288F0D866C;
        precomp_x[496] = 256'h3154137D779C25F14FF1FB88A6D0370B9E6AF48D88E7FC39C6417272EAA69B7C;
        precomp_x[497] = 256'hF8821E1FDFDF9FC81E3ACB3C1D1D7A65F710BE2D94A193550721CB9361549597;
        precomp_x[498] = 256'h8409463A521404A5A2D8AA90050E3AD8EC5D6FAF870333B06DD4F63E8354A655;
        precomp_x[499] = 256'h9680241112D370B56DA22EB535745D9E314380E568229E09F7241066003BC471;
        precomp_x[500] = 256'h9D1ABAEC9F5715A15C7628244170951E0F85E87F68CA5393D3F9FC3FA23A69C8;
        precomp_x[501] = 256'h1FB966918DB3AF46C37234B6A4B043719886D6A05859BA32F72742D6141F7AE6;
        precomp_x[502] = 256'h22D9E364B9274DAB098BCB23E0428E8A416D54F05A781281EE221DB69E1EC7B8;
        precomp_x[503] = 256'h625FA450AED083FB30166766D5874131ADB168C0247CBFF83987297BF873E45D;
        precomp_x[504] = 256'h24ACB1C19B6DFC25DEFB01C2E2681AE82DEACC0FF21AE8FF01F82F37A6A2147F;
        precomp_x[505] = 256'hD2856803A99D30D4F3A328E3BBF7DB3B6C6D1896BA5B339F33C1302CF75AB555;
        precomp_x[506] = 256'h80529E659D196884B15E95EF871E5FD88FB5298F3BC7831B50A0BC984CB5FE0A;
        precomp_x[507] = 256'h7F9199AA3B8201ED5D288E4949C432770E0BB316953F1DDED0674D7E8728E183;
        precomp_x[508] = 256'h7D32C88508E959F648C4674CDCCCB19129B4566D644D2FB76D0C89662C29ECBC;
        precomp_x[509] = 256'hF2B961C09291ECC8576CE67EBBD1BF011F1727FFAD9EB74CBF8819E32D1ABFBF;
        precomp_x[510] = 256'hD9A0C68995283291972D6A72897181B26B4AE3174E98A676F75BBFBF81BE876E;
        precomp_x[511] = 256'hC7A363246AEB7C8C991B2AA710ABDF5CFFF2991230B3A69FBE2DD4817C7C3E0A;
        precomp_y[0] = 256'h483ADA7726A3C4655DA4FBFC0E1108A8FD17B448A68554199C47D08FFB10D4B8;
        precomp_y[1] = 256'h388F7B0F632DE8140FE337E62A37F3566500A99934C2231B6CB9FD7584B8E672;
        precomp_y[2] = 256'hD8AC222636E5E3D6D4DBA9DDA6C9C426F788271BAB0D6840DCA87D3AA6AC62D6;
        precomp_y[3] = 256'h6AEBCA40BA255960A3178D6D861A54DBA813D0B813FDE7B5A5082628087264DA;
        precomp_y[4] = 256'hCC338921B0A7D9FD64380971763B61E9ADD888A4375F8E0F05CC262AC64F9C37;
        precomp_y[5] = 256'hD984A032EB6B5E190243DD56D7B7B365372DB1E2DFF9D6A8301D74C9C953C61B;
        precomp_y[6] = 256'h0AB0902E8D880A89758212EB65CDAF473A1A06DA521FA91F29B5CB52DB03ED81;
        precomp_y[7] = 256'h581E2872A86C72A683842EC228CC6DEFEA40AF2BD896D3A5C504DC9FF6A26B58;
        precomp_y[8] = 256'h4211AB0694635168E997B0EAD2A93DAECED1F4A04A95C0F6CFB199F69E56EB77;
        precomp_y[9] = 256'h85E89BC037945D93B343083B5A1C86131A01F60C50269763B570C854E5C09B7A;
        precomp_y[10] = 256'h321EB4075348F534D59C18259DDA3E1F4A1B3B2E71B1039C67BD3D8BCF81998C;
        precomp_y[11] = 256'h02DE1068295DD865B64569335BD5DD80181D70ECFC882648423BA76B532B7D67;
        precomp_y[12] = 256'h73016F7BF234AADE5D1AA71BDEA2B1FF3FC0DE2A887912FFE54A32CE97CB3402;
        precomp_y[13] = 256'hA69DCE4A7D6C98E8D4A1ACA87EF8D7003F83C230F3AFA726AB40E52290BE1C55;
        precomp_y[14] = 256'h2119A460CE326CDC76C45926C982FDAC0E106E861EDF61C5A039063F0E0E6482;
        precomp_y[15] = 256'hE022CF42C2BD4A708B3F5126F16A24AD8B33BA48D0423B6EFD5E6348100D8A82;
        precomp_y[16] = 256'hB9C398F186806F5D27561506E4557433A2CF15009E498AE7ADEE9D63D01B2396;
        precomp_y[17] = 256'h02972D2DE4F8D20681A78D93EC96FE23C26BFAE84FB14DB43B01E1E9056B8C49;
        precomp_y[18] = 256'h80FC06BD8CC5B01098088A1950EED0DB01AA132967AB472235F5642483B25EAF;
        precomp_y[19] = 256'h1C38303F1CC5C30F26E66BAD7FE72F70A65EED4CBE7024EB1AA01F56430BD57A;
        precomp_y[20] = 256'h0D0E3FA9ECA8726909559E0D79269046BDC59EA10C70CE2B02D499EC224DC7F7;
        precomp_y[21] = 256'hEECF41253136E5F99966F21881FD656EBC4345405C520DBC063465B521409933;
        precomp_y[22] = 256'h758F3F41AFD6ED428B3081B0512FD62A54C3F3AFBB5B6764B653052A12949C9A;
        precomp_y[23] = 256'h958EF42A7886B6400A08266E9BA1B37896C95330D97077CBBE8EB3C7671C60D6;
        precomp_y[24] = 256'hE0DEDC9B3B2F8DAD4DA1F32DEC2531DF9EB5FBEB0598E4FD1A117DBA703A3C37;
        precomp_y[25] = 256'h5ED430D78C296C3543114306DD8622D7C622E27C970A1DE31CB377B01AF7307E;
        precomp_y[26] = 256'hCEDABD9B82203F7E13D206FCDF4E33D92A6C53C26E5CCE26D6579962C4E31DF6;
        precomp_y[27] = 256'hCB474660EF35F5F2A41B643FA5E460575F4FA9B7962232A5C32F908318A04476;
        precomp_y[28] = 256'h4119B88753C15BD6A693B03FCDDBB45D5AC6BE74AB5F0EF44B0BE9475A7E4B40;
        precomp_y[29] = 256'h091B649609489D613D1D5E590F78E6D74ECFC061D57048BAD9E76F302C5B9C61;
        precomp_y[30] = 256'h0673FB86E5BDA30FB3CD0ED304EA49A023EE33D0197A695D0C5D98093C536683;
        precomp_y[31] = 256'h59C9E0BBA394E76F40C0AA58379A3CB6A5A2283993E90C4167002AF4920E37F5;
        precomp_y[32] = 256'h3B952D32C67CF77E2E17446E204180AB21FB8090895138B4A4A797F86E80888B;
        precomp_y[33] = 256'h55EB2DAFD84D6CCD5F862B785DC39D4AB157222720EF9DA217B8C45CF2BA2417;
        precomp_y[34] = 256'hEFAE9C8DBC14130661E8CEC030C89AD0C13C66C0D17A2905CDC706AB7399A868;
        precomp_y[35] = 256'hE38DA76DCD440621988D00BCF79AF25D5B29C094DB2A23146D003AFD41943E7A;
        precomp_y[36] = 256'hF98A3FD831EB2B749A93B0E6F35CFB40C8CD5AA667A15581BC2FEDED498FD9C6;
        precomp_y[37] = 256'h744B1152EACBE5E38DCC887980DA38B897584A65FA06CEDD2C924F97CBAC5996;
        precomp_y[38] = 256'hC534AD44175FBC300F4EA6CE648309A042CE739A7919798CD85E216C4A307F6E;
        precomp_y[39] = 256'hE13817B44EE14DE663BF4BC808341F326949E21A6A75C2570778419BDAF5733D;
        precomp_y[40] = 256'h30E93E864E669D82224B967C3020B8FA8D1E4E350B6CBCC537A48B57841163A2;
        precomp_y[41] = 256'hE491A42537F6E597D5D28A3224B1BC25DF9154EFBD2EF1D2CBBA2CAE5347D57E;
        precomp_y[42] = 256'h100B610EC4FFB4760D5C1FC133EF6F6B12507A051F04AC5760AFA5B29DB83437;
        precomp_y[43] = 256'hEF0AFBB2056205448E1652C48E8127FC6039E77C15C2378B7E7D15A0DE293311;
        precomp_y[44] = 256'h8B378A22D827278D89C5E9BE8F9508AE3C2AD46290358630AFB34DB04EEDE0A4;
        precomp_y[45] = 256'h68651CF9B6DA903E0914448C6CD9D4CA896878F5282BE4C8CC06E2A404078575;
        precomp_y[46] = 256'hF5435A2BD2BADF7D485A4D8B8DB9FCCE3E1EF8E0201E4578C54673BC1DC5EA1D;
        precomp_y[47] = 256'hD56EB30B69463E7234F5137B73B84177434800BACEBFC685FC37BBE9EFE4070D;
        precomp_y[48] = 256'hEDD77F50BCB5A3CAB2E90737309667F2641462A54070F3D519212D39C197A629;
        precomp_y[49] = 256'h0A855BABAD5CD60C88B430A69F53A1A7A38289154964799BE43D06D77D31DA06;
        precomp_y[50] = 256'h66DB656F87D1F04FFFD1F04788C06830871EC5A64FEEE685BD80F0B1286D8374;
        precomp_y[51] = 256'h09414685E97B1B5954BD46F730174136D57F1CEEB487443DC5321857BA73ABEE;
        precomp_y[52] = 256'h4CB95957E83D40B0F73AF4544CCCF6B1F4B08D3C07B27FB8D8C2962A400766D1;
        precomp_y[53] = 256'hFA77968128D9C92EE1010F337AD4717EFF15DB5ED3C049B3411E0315EAA4593B;
        precomp_y[54] = 256'h5F3032F5892156E39CCD3D7915B9E1DA2E6DAC9E6F26E961118D14B8462E1661;
        precomp_y[55] = 256'h8EC0BA238B96BEC0CBDDDCAE0AA442542EEE1FF50C986EA6B39847B3CC092FF6;
        precomp_y[56] = 256'h8DC2412AAFE3BE5C4C5F37E0ECC5F9F6A446989AF04C4E25EBAAC479EC1C8C1E;
        precomp_y[57] = 256'h5E4631150E62FB40D0E8C2A7CA5804A39D58186A50E497139626778E25B0674D;
        precomp_y[58] = 256'hF65F5D3E292C2E0819A528391C994624D784869D7E6EA67FB18041024EDC07DC;
        precomp_y[59] = 256'hF3E0319169EB9B85D5404795539A5E68FA1FBD583C064D2462B675F194A3DDB4;
        precomp_y[60] = 256'h42242A969283A5F339BA7F075E36BA2AF925CE30D767ED6E55F4B031880D562C;
        precomp_y[61] = 256'h204B5D6F84822C307E4B4A7140737AEC23FC63B65B35F86A10026DBD2D864E6B;
        precomp_y[62] = 256'h04F14351D0087EFA49D245B328984989D5CAF9450F34BFC0ED16E96B58FA9913;
        precomp_y[63] = 256'h073867F59C0659E81904F9A1C7543698E62562D6744C169CE7A36DE01A8D6154;
        precomp_y[64] = 256'h39F23F366809085BEEBFC71181313775A99C9AED7D8BA38B161384C746012865;
        precomp_y[65] = 256'hD2424B1B1ABE4EB8164227B085C9AA9456EA13493FD563E06FD51CF5694C78FC;
        precomp_y[66] = 256'hEAD12168595FE1BE99252129B6E56B3391F7AB1410CD1E0EF3DCDCABD2FDA224;
        precomp_y[67] = 256'h6FDCEF09F2F6D0A044E654AEF624136F503D459C3E89845858A47A9129CDD24E;
        precomp_y[68] = 256'h060660257DD11B3AA9C8ED618D24EDFF2306D320F1D03010E33A7D2057F3B3B6;
        precomp_y[69] = 256'h3D98A9CDD026DD43F39048F25A8847F4FCAFAD1895D7A633C6FED3C35E999511;
        precomp_y[70] = 256'h0B4C4FE99C775A606E2D8862179139FFDA61DC861C019E55CD2876EB2A27D84B;
        precomp_y[71] = 256'hAE434102EDDE0958EC4B19D917A6A28E6B72DA1834AFF0E650F049503A296CF2;
        precomp_y[72] = 256'hCF2174118C8B6D7A4B48F6D534CE5C79422C086A63460502B827CE62A326683C;
        precomp_y[73] = 256'h6FB8D5591B466F8FC63DB50F1C0F1C69013F996887B8244D2CDEC417AFEA8FA3;
        precomp_y[74] = 256'h322AF4908C7312B0CFBFE369F7A7B3CDB7D4494BC2823700CFD652188A3EA98D;
        precomp_y[75] = 256'h6749E67C029B85F52A034EAFD096836B2520818680E26AC8F3DFBCDB71749700;
        precomp_y[76] = 256'h2AEABE7E4531510116217F07BF4D07300DE97E4874F81F533420A72EEB0BD6A4;
        precomp_y[77] = 256'hB0EA558A113C30BEA60FC4775460C7901FF0B053D25CA2BDEEE98F1A4BE5D196;
        precomp_y[78] = 256'h998C74A8CD45AC01289D5833A7BEB4744FF536B01B257BE4C5767BEA93EA57A4;
        precomp_y[79] = 256'hB2284279995A34E2F9D4DE7396FC18B80F9B8B9FDD270F6661F79CA4C81BD257;
        precomp_y[80] = 256'hBDD46039FEED17881D1E0862DB347F8CF395B74FC4BCDC4E940B74E3AC1F1B13;
        precomp_y[81] = 256'h6F0A256BC5EFDF429A2FB6242F1A43A2D9B925BB4A4B3A26BB8E0F45EB596096;
        precomp_y[82] = 256'hC359D6923BB398F7FD4473E16FE1C28475B740DD098075E6C0E8649113DC3A38;
        precomp_y[83] = 256'h021AE7F4680E889BB130619E2C0F95A360CEB573C70603139862AFD617FA9B9F;
        precomp_y[84] = 256'h60EA7F61A353524D1C987F6ECEC92F086D565AB687870CB12689FF1E31C74448;
        precomp_y[85] = 256'h49B96715AB6878A79E78F07CE5680C5D6673051B4935BD897FEA824B77DC208A;
        precomp_y[86] = 256'h5CA560753BE2A12FC6DE6CAF2CB489565DB936156B9514E1BB5E83037E0FA2D4;
        precomp_y[87] = 256'h7571D74EE5E0FB92A7A8B33A07783341A5492144CC54BCC40A94473693606437;
        precomp_y[88] = 256'hBE52D107BCFA09D8BCB9736A828CFA7FAC8DB17BF7A76A2C42AD961409018CF7;
        precomp_y[89] = 256'h8FD64A14C06B589C26B947AE2BCF6BFA0149EF0BE14ED4D80F448A01C43B1C6D;
        precomp_y[90] = 256'h39E5C9925B5A54B07433A4F18C61726F8BB131C012CA542EB24A8AC07200682A;
        precomp_y[91] = 256'h62DFAF07A0F78FEB30E30D6295853CE189E127760AD6CF7FAE164E122A208D54;
        precomp_y[92] = 256'h25A748AB367979D98733C38A1FA1C2E7DC6CC07DB2D60A9AE7A76AAA49BD0F77;
        precomp_y[93] = 256'hECFB7056CF1DE042F9420BAB396793C0C390BDE74B4BBDFF16A83AE09A9A7517;
        precomp_y[94] = 256'hCD450EC335438986DFEFA10C57FEA9BCC521A0959B2D80BBF74B190DCA712D10;
        precomp_y[95] = 256'hF5C54754A8F71EE540B9B48728473E314F729AC5308B06938360990E2BFAD125;
        precomp_y[96] = 256'h6CB9A8876D9CB8520609AF3ADD26CD20A0A7CD8A9411131CE85F44100099223E;
        precomp_y[97] = 256'hFEF5A3C68059A6DEC5D624114BF1E91AAC2B9DA568D6ABEB2570D55646B8ADF1;
        precomp_y[98] = 256'h1ACB250F255DD61C43D94CCC670D0F58F49AE3FA15B96623E5430DA0AD6C62B2;
        precomp_y[99] = 256'h5F310D4B3C99B9EBB19F77D41C1DEE018CF0D34FD4191614003E945A1216E423;
        precomp_y[100] = 256'h438136D603E858A3A5C440C38ECCBADDC1D2942114E2EDDD4740D098CED1F0D8;
        precomp_y[101] = 256'hCDB559EEDC2D79F926BAF44FB84EA4D44BCF50FEE51D7CEB30E2E7F463036758;
        precomp_y[102] = 256'h0C3B997D050EE5D423EBAF66A6DB9F57B3180C902875679DE924B69D84A7B375;
        precomp_y[103] = 256'h6D89AD7BA4876B0B22C2CA280C682862F342C8591F1DAF5170E07BFD9CCAFA7D;
        precomp_y[104] = 256'hCA5EF7D4B231C94C3B15389A5F6311E9DAFF7BB67B103E9880EF4BFF637ACAEC;
        precomp_y[105] = 256'h09731141D81FC8F8084D37C6E7542006B3EE1B40D60DFE5362A5B132FD17DDC0;
        precomp_y[106] = 256'hEE1849F513DF71E32EFC3896EE28260C73BB80547AE2275BA497237794C8753C;
        precomp_y[107] = 256'hD3AA2ED71C9DD2247A62DF062736EB0BADDEA9E36122D2BE8641ABCB005CC4A4;
        precomp_y[108] = 256'hC4E1020916980A4DA5D01AC5E6AD330734EF0D7906631C4F2390426B2EDD791F;
        precomp_y[109] = 256'h67163E903236289F776F22C25FB8A3AFC1732F2B84B4E95DBDA47AE5A0852649;
        precomp_y[110] = 256'h0CD1BC7CB6CC407BB2F0CA647C718A730CF71872E7D0D2A53FA20EFCDFE61826;
        precomp_y[111] = 256'h299D21F9413F33B3EDF43B257004580B70DB57DA0B182259E09EECC69E0D38A5;
        precomp_y[112] = 256'hF9429E738B8E53B968E99016C059707782E14F4535359D582FC416910B3EEA87;
        precomp_y[113] = 256'h462F9BCE619898638499350113BBC9B10A878D35DA70740DC695A559EB88DB7B;
        precomp_y[114] = 256'h62188BC49D61E5428573D48A74E1C655B1C61090905682A0D5558ED72DCCB9BC;
        precomp_y[115] = 256'h7C10DFB164C3425F5C71A3F9D7992038F1065224F72BB9D1D902A6D13037B47C;
        precomp_y[116] = 256'hAB8C1E086D04E813744A655B2DF8D5F83B3CDC6FAA3088C1D3AEA1454E3A1D5F;
        precomp_y[117] = 256'h4CB04437F391ED73111A13CC1D4DD0DB1693465C2240480D8955E8592F27447A;
        precomp_y[118] = 256'hBD1AEB21AD22EBB22A10F0303417C6D964F8CDD7DF0ACA614B10DC14D125AC46;
        precomp_y[119] = 256'hBFEFACDB0E5D0FD7DF3A311A94DE062B26B80C61FBC97508B79992671EF7CA7F;
        precomp_y[120] = 256'h603C12DAF3D9862EF2B25FE1DE289AED24ED291E0EC6708703A5BD567F32ED03;
        precomp_y[121] = 256'hCC6157EF18C9C63CD6193D83631BBEA0093E0968942E8C33D5737FD790E0DB08;
        precomp_y[122] = 256'h553E04F6B018B4FA6C8F39E7F311D3176290D0E0F19CA73F17714D9977A22FF8;
        precomp_y[123] = 256'h0712FCDD1B9053F09003A3481FA7762E9FFD7C8EF35A38509E2FBF2629008373;
        precomp_y[124] = 256'hED8CC9D04B29EB877D270B4878DC43C19AEFD31F4EEE09EE7B47834C1FA4B1C3;
        precomp_y[125] = 256'h9852390A99507679FD0B86FD2B39A868D7EFC22151346E1A3CA4726586A6BED8;
        precomp_y[126] = 256'h9E994980D9917E22B76B061927FA04143D096CCC54963E6A5EBFA5F3F8E286C1;
        precomp_y[127] = 256'h4036EDC931A60AE889353F77FD53DE4A2708B26B6F5DA72AD3394119DAF408F9;
        precomp_y[128] = 256'h753C8B9F9754F18D87F21145D9E2936B5EE050B27BBD9681442C76E92FCF91E6;
        precomp_y[129] = 256'h86CA160D68F4D4E718B495B891D3B1B573B871A702B4CF6123ABD4483AA79C64;
        precomp_y[130] = 256'h8147CBF7B973FCC15B57B6A3CFAD6863EDD0F30E3C45B85DC300C513C247759D;
        precomp_y[131] = 256'h31B3CA455073BEA558ADBE56C27B470BAF949AE650213921DC287844F1A29574;
        precomp_y[132] = 256'h57FC24472225B23F5714626D8D67D56110BD3A60DD7A16870CBBB893F652F50F;
        precomp_y[133] = 256'h844ADB5CE7D10DE94617C73CA77040E4EE4E92E0156B3C70CC593FA494B33482;
        precomp_y[134] = 256'hD765466C6E556E352F77872225627D80A73538074B44FF27057AD22E2F2454A2;
        precomp_y[135] = 256'h77B1F0687CFCDBE8812605E50D8B752CDA811844236A4C4377F53C946E7BD648;
        precomp_y[136] = 256'hC16F60C7C11FC3C9EB27FA26A9035B669BFB77D21CEF371DDCE94E329222550C;
        precomp_y[137] = 256'hE1BCFE7FC8ED8AE95CF6C2437FDD94BFD742E8CAA6DE78114C25112A86988EFD;
        precomp_y[138] = 256'h8D6857C9D08EF7B4FD8883363D37BEE70FE8529F7173F58943FCAE81D2D0EA0E;
        precomp_y[139] = 256'hDDF1B9FE8744AD03F996BF6B96EC34962B601BD5ED952F7854F583888917BE80;
        precomp_y[140] = 256'h3F27E7E1834F1A61AF6F04DC61E7AE64716BC5E0A6B063B301D0E60E47298A9D;
        precomp_y[141] = 256'h50BC23F3926CD0C49F53FBB235EB1E890D579517F5BDC3AB2416DB785AAEDB3F;
        precomp_y[142] = 256'h6E6AEE6C9625370AF866C25C7CA5DD780527EFBCE7D8B3A39AB249309A185187;
        precomp_y[143] = 256'h986314EF75B68FB2827C2965041981395D699FCD81CF23CE7019BC4135174870;
        precomp_y[144] = 256'h4E31EA12AC607D075DE4B22DE1BE2C52E0A44D254728D2C544D2DDF9E3E469C0;
        precomp_y[145] = 256'h94264621A5960E0EE24C27926F16CAD2907F2636762E8D5A17E94AFD8E9D2BB0;
        precomp_y[146] = 256'h5B5853AB7EE5DE8D34E3D6BEB201094FFF8FBD1E0682F7F1EF87DDD65D7303C9;
        precomp_y[147] = 256'h496C944DD9875BA60A537EF96BF4C714A0AFFF24387D95E89B42337A33110753;
        precomp_y[148] = 256'hF2ECCAC775922B50899C979A02B3CC30B629E62E85693BA470F6EE381284C162;
        precomp_y[149] = 256'h44C757A542F4EA2EB39605D4268C2510AC685AABD77A8F5C4D95E23F4C2E9368;
        precomp_y[150] = 256'h7421A2207EE73299D46192FC93CA03DEC824ED8DE2F48367EC5383170A17FFFB;
        precomp_y[151] = 256'h7D16D654F0C2AFF0FC254DAD063761A26C8D4022EA85B8CC22F3EA1EF69961A9;
        precomp_y[152] = 256'h6C9ED1F1528B021593A39839340DDB530A2F2E365290C49824B035C673C9259D;
        precomp_y[153] = 256'h0E8BCBFE1F7F6E75D32E20499329765F02EFFC56A922F26860D4BC0AADD0E24D;
        precomp_y[154] = 256'h3E18941CC3C6D297CC9A32F695807B1C7DA8561DE4FDE71D4F9BBDB6E9BF3916;
        precomp_y[155] = 256'hF60547AB6E9C5FD3ECA6E349B85880C61FDAD0FC2F7AB155295CAAECB973C154;
        precomp_y[156] = 256'h29A835F6EF7FA1E5F6F37A80CF96CA9843762BB1B12A0DAEAE83234BD0B5CCD5;
        precomp_y[157] = 256'h5C7BCF8B57F114E0B73BCFB810F5C60D35DC99AE9DC7F0E2606CC1F728C2071E;
        precomp_y[158] = 256'hA286E222DFE10CFD9689EABA6A81F04489C86DB6869AA1B554A90F1E83778EEE;
        precomp_y[159] = 256'hC582DB1A3F0F22421913B2E951E98A78660B4C40AD08FD65528593BC18223188;
        precomp_y[160] = 256'hE3E77C41288F2602E722AF7F4B70E64DE4116FB9955B03B06EA8B19F7A20350D;
        precomp_y[161] = 256'hC9E33FAEBD8EBA426736C0C76F3DEABAEE2B59C50953FB43C2DCC5139E7C4BDC;
        precomp_y[162] = 256'hF5202CF5AAEEA58BF4F58C7EDF4417BE1B87FFDEE68E77F0D7E81ABE158E3A25;
        precomp_y[163] = 256'h61FE64CAB0952CAE3C574F282F74A87DC2A96316B7009F2E4E9C5FCC12285844;
        precomp_y[164] = 256'h5DCF9ABBA9625ED680B0F20FB1F047D593A0C61C539692538CDF6B034D730B58;
        precomp_y[165] = 256'h79A6BF4375F1469C4F5321C6C72FBBF4BA7CEC105675F437B5E013AD7B5D75D4;
        precomp_y[166] = 256'h7669BBD419A4D491F592A35B6AA3DFE45BD2FE7FD179C7781CD5F918D732F63D;
        precomp_y[167] = 256'h308ABC8DF271F75959B20C5C7FA62BAFBFC9CCBF49B946A954E5381C1728D1C7;
        precomp_y[168] = 256'h9EEA970BA856B2FAA3E82877CC84ED4F3DC0EFBA1E7C3BAA8B386FFC46E0AE7E;
        precomp_y[169] = 256'hA9FB1702100953B359B2E2688AE7FD33A30377DA47BFDA713E2D7D73DFB1030C;
        precomp_y[170] = 256'h22F6FE9D217495017FDB7F5B2F12FA57095F40E131714885C12A2EA16EDB6BE6;
        precomp_y[171] = 256'h737CECA2C0EF72278B90501CCB71B6715E5C31D4CD0478C118FE128795F1DD0C;
        precomp_y[172] = 256'h2AFC8D09B79176D8D003FD2A4F18D526403FFF272D47E7787376FEB7CBDDD8FD;
        precomp_y[173] = 256'hCB13C152FD511D91A9E0ED90AFA021A081F77F6D20CC1376E2195FFCF28FA758;
        precomp_y[174] = 256'h1AB4EABE5E09409D75CCA8922647F48DBD698A16D4F7CC8596DAF16940023A52;
        precomp_y[175] = 256'h95F9F4E9007E5B9FA48FA422A26AB982DC48A4D54D7123986E6D3AB974E88915;
        precomp_y[176] = 256'hDCE1BAE1D655BA517F5B5580997117570A77CD3BDD4B8E8E330E97791BC31DF0;
        precomp_y[177] = 256'hCC3636A03FDDDDFABED88DAAB081F3591C48D2CA71BA34FCF6989F4AF7625D8E;
        precomp_y[178] = 256'h329CF0497E15EEC7B8EAFC4A0B8A7D1CD8B632038D4AEF81974CF9844611A32D;
        precomp_y[179] = 256'h8C6F81BE3FAFA5EEC8296F928AC7919DC4D88C9A59442274D0531B7BF7E48E78;
        precomp_y[180] = 256'h7F42C0962FEB2F73B2B0965A1F359A6ADE49D768A2CE6B07B5ACB92B73E05583;
        precomp_y[181] = 256'hF649BE278CAD976420742CE382DCE3A1420E372EF1B25B2759A8ED387282765E;
        precomp_y[182] = 256'hD596ADF0E8692A06BC6284BF0299BEF685E2A171585AA1324B9A05B50CE815B7;
        precomp_y[183] = 256'hE077184B4AE8F7056C10DD9EF541689D143F6871789E1801DEAEFC1D527A8FB4;
        precomp_y[184] = 256'hEB4C98489093D573A295407E1D6FC48A787120CEB3D3DCFBB40634E0E75E221D;
        precomp_y[185] = 256'hEA75B9B25D717861D1AF1C019C372941C8968B90EF134F9F323215E1BB0B2155;
        precomp_y[186] = 256'h669985206EDF4AC6F39BE21F20C98824210E204CE44998095DE355371641218C;
        precomp_y[187] = 256'h70B0123774AF550E68E68E5F65CA6E9808846E03CF39AF778511BE82BC32FEFE;
        precomp_y[188] = 256'hE115B14BEF4695CFFB85BDF98BA3985CBD5E5B8983E053907C36F9CE8B75D41D;
        precomp_y[189] = 256'hE9D9DBFE8CF5F5CCA855D6CCBD11F48060FAFA8DAD6BD3E9C86DF5CEB0FA5270;
        precomp_y[190] = 256'hE4177CE1C3CD6AC778925BD67E72CB77D1925B91D06A7F1698411A4786393FB0;
        precomp_y[191] = 256'h954A5FD857BA3ACF2D4B1F41E8E1F2CD1F21C4B96899781B742A49D2E61ED18B;
        precomp_y[192] = 256'h2D5D2FB1F0C308553B1FE249298B2059259D3D49D4D7071ADCE4BCC5DC937193;
        precomp_y[193] = 256'h9BD0178E381895692217267B7407E98727FCAEDA12D8CF5449EB5472D554E0FF;
        precomp_y[194] = 256'h618BD6B0D25CA70DF08B76929336E421691B09730F2F5A052E7ADC173584427B;
        precomp_y[195] = 256'h07A981F0C21862A853B4F895DC62482C530ED7385E5D1E330CFB9D0FE879992C;
        precomp_y[196] = 256'hADB23BCDB3D069C5E83BE30B2469B0680B2A81B7B667E934233B75EFB5753F28;
        precomp_y[197] = 256'hD8003C9EE3C842F5EDE375A8A7768DB4803ECF119B7B37DECEA15631B4E8DBCA;
        precomp_y[198] = 256'h211557489FA93B883E5BEA50DA005C5368E21A0C41BC83D9145C13E1370D26D0;
        precomp_y[199] = 256'hABB1D9F874637668E214EFBAFBF529D312FF023BC1D5723E585404366834F189;
        precomp_y[200] = 256'h5B5930F12E9C40BCB3393A895C2D64576A3ABD23B7291B99C965C33DEF60A55C;
        precomp_y[201] = 256'h5246A8190BBFB2915F82ED5650796F505CED5C2587347D57A873CEAF3D997E7A;
        precomp_y[202] = 256'h3C83145DAD9F87487B97E7464850ED02D71DBD04093281A13D2127766A791EE2;
        precomp_y[203] = 256'h6CE693B64A37C6727E141041AB9A0D589AB9C303A5AC3D3EC89B6F279E79827C;
        precomp_y[204] = 256'hF602C3428593A9A8D671D1BC7C1D88340FE9F5F52E6A7F0FBB8701464E6F4838;
        precomp_y[205] = 256'hB8F7C3B220701320F20CA036761D3E56BF94A7009A919F1A3EA0CB81B74424A6;
        precomp_y[206] = 256'hAFB6A74D9849454EDD7F703A5C6616D143F9CBCC9A9A5D6F6A7B5D1F9D9FCAFF;
        precomp_y[207] = 256'hDA7D67CBC1EDE9D4FEDD5DCDC96B04F9A3561BA02581B055EAA144EB4217DACA;
        precomp_y[208] = 256'h160E1C1C13342FD459D4F9898AE632B842B8947913733B89384FC1042D30BF01;
        precomp_y[209] = 256'h87092DCBB9C3D254E3B055FF3A76EC0564C4A7C57FB1783CEFDC40FC10B751F0;
        precomp_y[210] = 256'hFE49A6A8B5E46BF1EF679714DABD590EA831D46B8EE94EB613132BA37855FABB;
        precomp_y[211] = 256'h4521954EFCC98263DF2F14E0E6E6B47AF6B83F0BBC20722C15445F87E05F4513;
        precomp_y[212] = 256'hCD15ABBCD744D4850D5E401F1F89A5DF122F37B4E362B4CEE3E53B1C00110BF3;
        precomp_y[213] = 256'hCFD4D36BEB2E11F241FD0F367A0737AD303E915FF247F131368CA50918E00957;
        precomp_y[214] = 256'h72EA16B532A7336D3332400B303C0236B6A1294D88CE7FE915571284D1F7C189;
        precomp_y[215] = 256'hD5E6268B30952422BE59FE0EFE7BA2E703215994827A46C2F2972B26153CF7AE;
        precomp_y[216] = 256'hB8241453ABC44C57DDAD6FF386D416F43E258A390C6F88379F80472B943F32B9;
        precomp_y[217] = 256'hC1FDAC5AEF4C6F0FFCB8E1C5C4417C713E3D5F07146DAA1AAAF2E7FEE70C4914;
        precomp_y[218] = 256'hFD5A31976FAD6AEEC304752CC3EBBC511F3695B09A737FA30AF42CC6EFD684CC;
        precomp_y[219] = 256'h563651760897632F8DDE31677A24F55834C5C9A55C1CBF36FD8B44803C9C6C81;
        precomp_y[220] = 256'hB5CE31605D6DD9C622CAE425CCD28912C4439820C06950CD4C86D9B453ABD7ED;
        precomp_y[221] = 256'h933D348378A71F443788194AAFC545E7F53E37A6F779F96E8FA14CCDEDE3B4EB;
        precomp_y[222] = 256'h2A7D3701A8724B12BD7C4830224AC083CBEA83D0543B541480BA8C8AE7731232;
        precomp_y[223] = 256'hEA90F8AAE214EE16ED608A72366998994E311DC7780EF885B29290C3823C470E;
        precomp_y[224] = 256'hCB7571C4071C552765BD289EA3CF3F38796DA2B12C953D0B8705125C4861D598;
        precomp_y[225] = 256'h7BBBB198EB39973B76D87F8194D45150A66D4F3B128A40BEC989A405AD7C287B;
        precomp_y[226] = 256'hA2F2F02A8272DE6E3DC8B39508959AD251B6D3D004C8195259A501E28FF7892A;
        precomp_y[227] = 256'h8613BB848398681D66F1E75D5B6EF44FD827B6290F4956A441D8F503DD32B289;
        precomp_y[228] = 256'h838E779334AA6FE6CAE90A62D359C339187B403215D97CDA4E62724AA5A50306;
        precomp_y[229] = 256'h01FCABF21E19CE68EE12A3D284BD1304010FA5F5D45F9C15D4070243A8433047;
        precomp_y[230] = 256'hE15723EB0E0BDBE6D6F28D6DA0443C634851F5B4C551BEC69F9196A00969ED71;
        precomp_y[231] = 256'hFFB0E211C79FBB7978BD4E53A05A267FF1E32C34D6287DEE64576D31AB959AB2;
        precomp_y[232] = 256'hF6A9186FF147B9B5FFC844B2EC0E255A1AE5537D75624288CE8421F87E94E1A4;
        precomp_y[233] = 256'h8791C0007C09C94DB328034B88C5BBBC113335366679EB099A5E75B583BC2C2A;
        precomp_y[234] = 256'h4B985B13C54990267FF564D2D4649C6F7E8FDBE1BA101D941C034E1464877B20;
        precomp_y[235] = 256'h31CE61A87834F52EFCF8703F93696F425813015563CA5D9CE92D8FC281135B0D;
        precomp_y[236] = 256'hBEA2A060505C13BC317CA083C5A8B85C9EAD5F6E1AC23FBEAC7CECEA9251C791;
        precomp_y[237] = 256'h74962C3FED9A6E9C896635EA855323B608850091F84DEE333CDFF8D0D2827928;
        precomp_y[238] = 256'h1CBCF83EA363E0D93E6ECC328653BA7AA165C526765B09F0696B0D61F122DB3A;
        precomp_y[239] = 256'hD10B5A637AB546BFCC610E2D1C3D61F461B0A806E7BA29C73D3DE909E9FAE659;
        precomp_y[240] = 256'h7B148EF273E1B131341AD4779342C7BC7B945A2CB52C448E4BB5FD503CEA1A19;
        precomp_y[241] = 256'h5847F4E06C6530335E29EA94389EE3E6D916314A60126028650AB9E0BFCFBBA7;
        precomp_y[242] = 256'h2CBFAD4D16C0702186611EEC408082FBFB2E9898141A52481C59E44ECD0676FF;
        precomp_y[243] = 256'h328E831D2F2B162C4ABE1644BB54CC8518DB178C5B6AE97E5E85110C7D7FDF1D;
        precomp_y[244] = 256'h627EEA93C6C9B53F9455941440A8B1006EBA68D46C922B6A1521F3946DD15E4E;
        precomp_y[245] = 256'h195A6A65D3790BEC716429863BCEF432E38242FC9F565DBBE159BC42F5740C69;
        precomp_y[246] = 256'h177C3A61682363ABBF281615D59F06FF5F87644C84D670E9A6C56AC1B611509B;
        precomp_y[247] = 256'h2D1A0B9C8EABA06543204DF148EB161825443EFA80F8AFF3D49B6626C5955AC8;
        precomp_y[248] = 256'h549B18C310FEAEA10225FADE934112D34058101D74F005381B82796AD0461736;
        precomp_y[249] = 256'hE95E050881AF550D09221F5AE95410316367D24BD545BDCB434E7638ACB46DBD;
        precomp_y[250] = 256'h62F637C67D8863748F1E2E26865118B999285B8755F25512C968B4FE49B8C971;
        precomp_y[251] = 256'hA0CBC0165E32171C8184265EAC7E0147206349D541035A94F56EFC49DCD7AB93;
        precomp_y[252] = 256'hA532D00D35013F859F4041D3AA231F2B9FC499670E0E2F824D5051F9E7F0C626;
        precomp_y[253] = 256'h92C20846CFDF1E8F3FE5BCAA06BDEDC39926833A3F40D28F23A8F952D8D18DDE;
        precomp_y[254] = 256'h1F023F2FA2BBECE703DBA14C124095CBFDC4F92F00281A148304A412C16ECAE6;
        precomp_y[255] = 256'h2DC6CAE5CAC2D88783DCA0E503C798F8FE067BCF5FC2975113756CF7EF4E5F1B;
        precomp_y[256] = 256'hB1DA863581531A1FBFB38A4E419FA1FECA8D55A83DDBCB98DA19D5CFFB7DA472;
        precomp_y[257] = 256'h4293260FE8AF6792A20B115EAA8376389094298B21D9DE16CF20E0C57A46089A;
        precomp_y[258] = 256'h5FC4756530E9B095F8B796431E745B991525BD4C04764E8EE8AF4B969BD6DDF6;
        precomp_y[259] = 256'hE1E79263A5BBBA8ACD78C92CFAECCD3AB84944D3785C07813763BF1ACE96C9DA;
        precomp_y[260] = 256'hF82B7D0E08EF9620E48C9F1353A72A95A9E11A3C1678CF10576E639BB1A7D04E;
        precomp_y[261] = 256'h86389E98E3C823C9E1B5384FFCE428C362E365797202FDBADC3D8C49395E7473;
        precomp_y[262] = 256'hF1D6314B661D1F8D8531D57B9470FB53D1509B2DA626A0FC4CAFC941B668BE84;
        precomp_y[263] = 256'hC296E64632F97DD5BA3B7012EAD44B6F324FCFD2F35F8B248E58FE68888BD453;
        precomp_y[264] = 256'hAC3B7747DE38C00F145FDB741482BB52324127CD2979EE12D4A9E689B9F8E778;
        precomp_y[265] = 256'h2DD3A45B94AAFE0753061CAA00A28560BD952B0B02F63F1396F42FB78E02FEF3;
        precomp_y[266] = 256'h00A873D9E70FD14AC2777A8FB5A02922BAE3A31A14938E69CB535355DE1EFADD;
        precomp_y[267] = 256'h14FE2225BF2BA0CC28C1C409E9849C4AD8ADF79263869B6854A28AE9631941FB;
        precomp_y[268] = 256'h24566B2455BC454AE7B378CCA0E57B6A8B821C8CA76FB858BB616E178907BE5A;
        precomp_y[269] = 256'h2A1125A2AC9968702BA22B5AD230C40E4E5C7E55D8BA6BA15E54D3CC7B72F3CC;
        precomp_y[270] = 256'h671FE16F00A65128591249E20B5070BF2A689E2BDD6C57DC18E5309AB6A40D0C;
        precomp_y[271] = 256'hAEC5402A54517B4C1F344D14B1943E69D7541F10C45BD4832B02B059499A6CC1;
        precomp_y[272] = 256'h5CBBD1861F80A4BD3D58262DEBC58FFD1D278FB3B4D7FEC6208F628677845CDC;
        precomp_y[273] = 256'h7EF486C50BF23BFBFC6DC15A41C0673FA9D003E6E1D09A8E4BFFEE9DAE2021E0;
        precomp_y[274] = 256'hE1F25BB21662B16D6D28A629AD84385A43DF566C52924BFD11854A78B70C22F5;
        precomp_y[275] = 256'h2AFFE855388660D827671E89C82832B225FA2C9B29D559E237AF565CB4DC99C3;
        precomp_y[276] = 256'hEA69F7945C6BABFF23400FD4A95D6833ABB27269887C372D8A6A45CAB25651AF;
        precomp_y[277] = 256'h6FF970A217BF47F80DA0AEABCB490E3B46C6DF3F69F9E93C3C4DD94AE7C05345;
        precomp_y[278] = 256'h9D6A55149867725A607A1C96EB03120CA497093934E0CF4A1631A63ABAC5DDB3;
        precomp_y[279] = 256'hF8A337C43181E3D569EC99D7F2BC4770CB6703A863FBD95B41FDB07CB697B447;
        precomp_y[280] = 256'h1B26ED76964DCF1B3F7FE6F32E6DB7E68E8FF4EE48FE63AF48FFD33BCD1645FE;
        precomp_y[281] = 256'h87640B41DBD99D16578A3D06D23D40888768A4E6DCF83E7B5B9D91335EB43D32;
        precomp_y[282] = 256'hFFED15017298FB9A78EB7BDF1430AC0482BAE82EA7197ADB50BCC1E1FC217B2E;
        precomp_y[283] = 256'hA9F8939B52AC53E35ED4771D8E47065C0D7F2805A7E5475C37353DDF182F4A65;
        precomp_y[284] = 256'h175D9B701C652EBF46B99F1F6E66C4A69B840019A48B1AC4878B386C03B7F81E;
        precomp_y[285] = 256'h1D457C0FA29D4C3FE65DED191127016DD40ADA90CBB0D8DEC2AF4BF820CC91DC;
        precomp_y[286] = 256'h7BC6B47090A7AFDBFC63905DDF69849973E1E4E2AF74F12663EAE8A4F4722D49;
        precomp_y[287] = 256'h7350EBAAF2CCF3C8F940CC14151C23C2BC33CB736552815692648F6B628E3FC8;
        precomp_y[288] = 256'h2E6E8B6BD83B7F5B1DC8E83BEDB3B23A80D9FF082029831A453050162BECE448;
        precomp_y[289] = 256'hC49C2A0095AEEE5B8DEB5E8CDB4D21E4CF0F31731AF2FAC525C534C234FFB328;
        precomp_y[290] = 256'hA0B67B7EBE8F59B3C25D546E03DC304DD22A6A64615BCFB925B685E318D43468;
        precomp_y[291] = 256'h2F51194352D07E517B7841F58EDA5225229A7E289A453AEB5E70110E12668436;
        precomp_y[292] = 256'h823FA47FA7B0B50C907056DC73E04574003F68A75A4C85668AB5F5B15657510B;
        precomp_y[293] = 256'h8DF4C9FAC94829EEFB0E7F521020B5B04F05F4D5839C86874E893E7D08AD92A3;
        precomp_y[294] = 256'hA030E8B6AC4E37A7DF01054AEA23A78E1BB7A22EF26052A3A034ECBCBC35ABDE;
        precomp_y[295] = 256'hCA18161D70360966CA381EA3F760B2FE28B040C7EBC82AF9BEA27BA6F4DFE8ED;
        precomp_y[296] = 256'hAEB27D0BEDF61FAC99528A9FF060D1F2376626B0BC807A19561C2E4FE8B49F65;
        precomp_y[297] = 256'h57D93436B354963C5891ABE3825D89B4D17685BCC9632E7EFE85DED75823C921;
        precomp_y[298] = 256'h13DAEFA0B2E2E09D36F472F229B5F7D158A18F63AC3DC4D6D62CC7D7EC0EF826;
        precomp_y[299] = 256'h867553EC17D2FD95B895EEDE15DA569ECBB3F25AE5F334A2B20660DFDF062383;
        precomp_y[300] = 256'hD5A7A1159900F90C879B1A3013945D8C5453BF1C07E5E33D6F8FAEAE439734EB;
        precomp_y[301] = 256'hDEBDA8597117EDE0DCC0ECC54EC1A494B3BBEE3495DB2B1EEBAA1DB92FC17C6F;
        precomp_y[302] = 256'h8BF48868E405D5332ADC0EC9049BC7CF1487E5543A043200717865218A39CC9D;
        precomp_y[303] = 256'h0D17E64ADD534A6EFDD0AF26B4494339F76B3C1B126397F9A2BEBA76EAF902AC;
        precomp_y[304] = 256'h7D9F38D474B5A22E72949F7FE2CEFB349A8FE1FBC16B8DDA11F162DE30E50F5B;
        precomp_y[305] = 256'h9BBBA8DD7C49204A9EDC4B91E38E4973FA61DE1CEDA6AD61603D97157F0B099D;
        precomp_y[306] = 256'hC26112CC006DCA2AFA52684FC9ED22D32F067891D5BAC2C02BB86E3B9411C61E;
        precomp_y[307] = 256'hB4EA854693FDE01CFB903A3118BB61F5C5047B94705A714D5B586D47A0142704;
        precomp_y[308] = 256'hDEB56AA5D45031EAFC411FECE09A964614664989FD4F40D779C0298198BBAB48;
        precomp_y[309] = 256'h2DAF9F3CEC44034FC8A71EE0EE76BD77AC6FDC9EFA042A2F6CAF9C5EFD130B97;
        precomp_y[310] = 256'h6BD0FD11F9E2DB7365F21DD134CB29F60FEF4D7FB419ABEFEAFE15A420DDB152;
        precomp_y[311] = 256'h7EA2FB40D460ADFFC9E25C530A65C508E77E6E76E2E435C2150C870A7600C823;
        precomp_y[312] = 256'h16E0958968066E52C873D6EFE549D3AA83D30BD6A1D730D368AA1AD232233145;
        precomp_y[313] = 256'h7EEACC27B2297FB563D691FA36DC650AF66FD3E66FE5E6379959D46E2D4BDDFA;
        precomp_y[314] = 256'h77593CC07E9D5E5E688A7B330BF54A01703CC9B7A0485E6D907515BB11A13FEF;
        precomp_y[315] = 256'hAD899E2250F6A8E8CE29B22583AD87552A6E6AB89061D33B6629FBFC52C0A241;
        precomp_y[316] = 256'h17E44EEB473F75BACFFAE683C8EA0299E19351807257803EF9963AD3D0989CE9;
        precomp_y[317] = 256'h7C55E76E8756796C143F64E7E40A402BEB537BE40F1F5322E59D2BE282776875;
        precomp_y[318] = 256'h782253186671273DA7B0B884E72E9BEE2B048C459430D2CA7C398AAA9FD9E2BC;
        precomp_y[319] = 256'h1759DB6388AED233CE0C5B47EC9DCB8876740928E12FE9D0D08EB7592D3F1990;
        precomp_y[320] = 256'h634C97ED0644A68FE1F1DA1F190CF9202B2DC810446B78EA9CD276843C76AAFD;
        precomp_y[321] = 256'h3A14266ABA263297FC6AB00A8403565DC9390B48EBFFCB6111B5E8EFC8F87182;
        precomp_y[322] = 256'hE4E6593A8E1AE842CA7F4EAED8CCCAA28A35F8DCCB8549BA2367FAF55F6C29C6;
        precomp_y[323] = 256'hFCA2C6BC4076C8EBA0978B9A2B0158C4338905142809461938413FE6C020385F;
        precomp_y[324] = 256'h007629F5AA367F51A29EBAF1235CF267F8016A6C88DFCD9B82D36904C949EAE2;
        precomp_y[325] = 256'h4F76B9FD24339C38C88C4217387B016DE4AE08FE67182D3982A45BB4E82BC60F;
        precomp_y[326] = 256'h9674AE58FE947C6D34C637252058C88C91B437DD98DA58B20EFD7E8D1615B9E5;
        precomp_y[327] = 256'h04C254541A5137425F75E515C04F1C73D11D50479C76B09BCE23C13ED1813251;
        precomp_y[328] = 256'hEC68E71C2E94E4904194753FD7484CA1940EAE5169831876877B9CE72D0B9DB1;
        precomp_y[329] = 256'h2915A9C5B770C86CEDD327493F698C176371F6A14CAC5A2273A3C6481B237FEF;
        precomp_y[330] = 256'hD3E6F8F16191DB06BE2274D15668589548E6925354F41114F43B5ED1013690C5;
        precomp_y[331] = 256'h608DFC157E3C23F44AA0FD883D02D2933C83EDCF066EA57F9167B7128D03DA21;
        precomp_y[332] = 256'h704967DF93FB862B3D38B18F4C6818AB6621C7D080D92CDD1F0092C0D7847903;
        precomp_y[333] = 256'hBF3B808EFE6B7EFB771853E56FBBA6E8B3B21FEF00706BD4274CC058B6FAE474;
        precomp_y[334] = 256'h9A424F366D3A79BE55BB5E9A283BE1E0163BFE221BC65E5E0318F0DE304D9AE7;
        precomp_y[335] = 256'h0CB478E6DFF8B9AA3AD06C6E8FC7E35A39BF6EC3787977BFD40F3159BF169E01;
        precomp_y[336] = 256'h032E3CDAEF60E55B0A9E36E6CD287737196C5AF8120C47B2F79D24929979263A;
        precomp_y[337] = 256'h2C396C5044A4953AB22A2D2247769741C5EDA54AD9C9AC97D6486B5F126DAC3E;
        precomp_y[338] = 256'h26D1D41225A1B5832DD53B9C56A6A8E8371DD19F31462DD9B2AEFE3E70412554;
        precomp_y[339] = 256'h40DEE344FC6F5C72C18B1603E149949CA0CFB31BB8B91B09C3CBABB0C6A5BFF0;
        precomp_y[340] = 256'h882E3A6DCACC1E928A3C1A6185F2BCF15E364F7A1EEEAAEA1C0AF593CF86185B;
        precomp_y[341] = 256'h72F61AE527B5C82E4AFA896655D9289D29931C1BF0D36C09FE4213C527848CBA;
        precomp_y[342] = 256'h0C3142CA54BCF2AE8B05DFB94E40F4BA7D3662F30774E61655C7515A87DDC5D5;
        precomp_y[343] = 256'hDAAE2D02041CABB20191B5BEC17E7E88957BFCD766DF1226A183064E3C4393A6;
        precomp_y[344] = 256'h98C35F7D69E5D98B920FFAFA6D15D3492D75FCB981CA50225AC7FF32618B1A20;
        precomp_y[345] = 256'h7175462EBE0F5EC007872B55356F2498976196BCEDBE021E08081EBDB2636298;
        precomp_y[346] = 256'h6E97EC27DD7D614DC1ED4FD8FDF6AA7008DCC3EBBE288831A9888166066333B2;
        precomp_y[347] = 256'hDADD16E764775BD5CA5C5F5135843556D7608230AAFF41254D4EAB381D28D2C0;
        precomp_y[348] = 256'h6EE1E84A77C6AB78A2CDA1B32FBDFE2E51D66843271D15C73F8E1A821E4C23A2;
        precomp_y[349] = 256'h092E7A5718EB0751C99254F4DDB5C278E17A417B21793339119A146DBBE3E0D3;
        precomp_y[350] = 256'hBAB4B2BA41BA4D53DF512E7632200BDC011D8583F2CEB5BDA8B7EB145CCC01FE;
        precomp_y[351] = 256'h3DDD27AFCD18049A3B01D0437761E4EA652FBD91115C470AE4C7BD4051EE73D2;
        precomp_y[352] = 256'h05DC9D46E5F6D94D48AF2EFC02F197A2F729F1D7335FA5690524D37C4ACD58C4;
        precomp_y[353] = 256'hB2683BF13FA8F7FCBE302823DFBC91538D902791D5D6DDE1D2805F370A0C08DB;
        precomp_y[354] = 256'hBAA8244C584FD05F2655E36BE2E5C459207D30EFDCDB229470B343339D16FF8F;
        precomp_y[355] = 256'h686FC317995446C4429452161A96595AA233B100E5F8BBC07199022944630BCD;
        precomp_y[356] = 256'h8961C913562385CA990593A377111A5D1DC6762BB1A928A66EBB304B8A24A701;
        precomp_y[357] = 256'h9CC24205ECF2708C357EDB54308CE45211F7DC0398FB48DB4982D33714C93046;
        precomp_y[358] = 256'hF65735B9708338C9ACC9CBA14B491B8AFB683058266A483D4987CDD389CCD0B4;
        precomp_y[359] = 256'h35039E3F8201E904E5378D032BD8B76626D9F0CE4425D2CEE7BBD24FB8725089;
        precomp_y[360] = 256'h58C58ECB7727A920B47A7E78E1E51D11E427D7E4465429BDA01F4650A4C102BB;
        precomp_y[361] = 256'hC2DEBC8958C3F60BD4C7B072D475A7D5C1EA784BC3E532BB72C0249009A42D65;
        precomp_y[362] = 256'hD389D64BB30BA9EB6CE80335CBE8F7DDB1EF3016A8B746602196B724D115605C;
        precomp_y[363] = 256'h49DB20A4D82397E56318640A6B605E9637D38961A58AE3DBFAC2FC11BBD11242;
        precomp_y[364] = 256'h8FF7E57CE79A08831FE8A9729249376407472B7761B055FA37105D18B51DF131;
        precomp_y[365] = 256'hBDEEEB418D2C4DC582547F6591C9721934778F5E0D25EFF494E243EDA6D34DA7;
        precomp_y[366] = 256'hAA23D2A47D6B717E55D7C6B65D9C46C68F2DB41CBA66960B4B4BF93F5FC88CB0;
        precomp_y[367] = 256'hCB079061353319B3A1669D59295BDBE218927D06CCB1290E4840CC16911A61D0;
        precomp_y[368] = 256'h2BFF7386527D6B5C2C595F80E08B4D2023BB8DFBF294DA12B54F8B14077281D0;
        precomp_y[369] = 256'h15BFD3BED3756AC6F2F1F9E60F254C9B2B1537171B2650816A2CC21B78B4DCF2;
        precomp_y[370] = 256'hC0111EDD3B4D28C4EDD264B8DC2BD0E320834DC7BDA82DD0827133C57F8CF73B;
        precomp_y[371] = 256'h9AFB5A57D71369C728DB308FB8B07DA0B91F954DB182EADB126B1FFFDDB673DA;
        precomp_y[372] = 256'hE7C99F66C49C8674A6C1B94B4B9640195E645CA7B3D2E0040AD8DC73F647CA5F;
        precomp_y[373] = 256'hA906AEECF901A3767D721F45DA53E3423BC0A779870E33C3D10F64266A2C8865;
        precomp_y[374] = 256'h403804C94339AE272BAFD894E63A4EB4690C1B4C9289DB00761E9B3A1D483F65;
        precomp_y[375] = 256'hB5C5FDDB332BFB59835E9A234AFA45435728DFAA7DCFCA3EA3C57DEBE849B336;
        precomp_y[376] = 256'h587B2E1F2E8EB9CB37AA6977870214EC818FB71C1035EECA91D53E68150CE67B;
        precomp_y[377] = 256'hCEE7991016A28462AA9DA7C00F67B4C7E8B3DD380F4B22039D05115AAC661DB8;
        precomp_y[378] = 256'h25952DAC4E1B50359B47E9B552852D1F300FDE75A6BD532F09FD56AF2A0AB333;
        precomp_y[379] = 256'hF527B8FD92234151BA11F24F7BD5DFED6EBD03E3A5048C6E8F2D52317201BAFE;
        precomp_y[380] = 256'h275CC76486C86A900F597DD67092ECFF5382C7B733939CA1D1F3218D6F0B594B;
        precomp_y[381] = 256'hB5EBE8FFB30DE5BDA532604416ABBAE14FF9198EB491794AC4500031947A985D;
        precomp_y[382] = 256'h2475618998BB414D4A534C6BE300297BAADF4FFCB10E67954EA36E252CF3CAC0;
        precomp_y[383] = 256'hD9FC5AB2CD619D4AC66C1CD2251504CCCDA34A7686C5661A960A00F8E4AA7E66;
        precomp_y[384] = 256'hD7D8DF98442060E00F17A363579C6600360B51242774E2DFC8D4B7871E1874E7;
        precomp_y[385] = 256'h470DCFD7B0C8C2ED63A28074A505573B42F509206B0AE57727A8B7967A0F42B1;
        precomp_y[386] = 256'h2F78934602A636A99BA2A1D232829F4139B579670BB26D0C898798BB6521D439;
        precomp_y[387] = 256'h326409B070550E9758F536987936A54AB701F7B678A7D10FEBB511A6C18CC917;
        precomp_y[388] = 256'h1B251CA52AF897AC4C08DF48CE3D1607D3B31B2C2DCD7F7A59A95B07774C4D83;
        precomp_y[389] = 256'hF4FB60B074419630FBAF5B53717B2A6F5CC2D98F1D29481B77B1F9F384175729;
        precomp_y[390] = 256'h635A39530046FBBF903DC729D3E3B52B43EEBDC53748ED833C95EAF71B75790F;
        precomp_y[391] = 256'h4983C08BF2D81C52D3B3A202E0C6DDB932A43A45C4B95F82C8C106425A783B52;
        precomp_y[392] = 256'h561EE03245CC3066968853F751FA36BE0CB50740A5951E87CF77EF20CB27E110;
        precomp_y[393] = 256'hF2B23CFF05EBDC8C0558DB8C1C311A94E9D8F63AD1CF4AF4C21C2349A6E57C4C;
        precomp_y[394] = 256'h950499C019719DAE0FDA04248D851E52CF9D66EEB211D89A77BE40DE22B6C89D;
        precomp_y[395] = 256'h9B03C7579704E839C8EEC7D0F063C4FDD0AA7BA05AD75254984B1703AE69A3D6;
        precomp_y[396] = 256'h26EF6B3D7B037663979333FE056BC33ACA54A3DD78C9244D79EF5426F2B69A02;
        precomp_y[397] = 256'h8BCC1D05FB880EC78762D8F3F5AFEFE8F4345BD836397D23BEFDF446498511C3;
        precomp_y[398] = 256'h2E6A15E11F77633530FB2CDB788AAA9883105DA307E28C0A8FAD503EB9779DF2;
        precomp_y[399] = 256'h08F7ABF1103E92F55DCB1DDE746DF10DA86BFB8D2776A0F01D07142DC9BCA443;
        precomp_y[400] = 256'h82EEB8A10F0B966FBBC3858A3878F969A853E2BBE1B60C4EE13EFF850D2D2CA7;
        precomp_y[401] = 256'h28F9D653C4042478831CCFE7BEC866635E0D32EDF6DB4F5425669A91D1DC0193;
        precomp_y[402] = 256'h05ABC582274876D63DCE366AFBB1D80A2286DC2ADC0C078F1424D45E026666B3;
        precomp_y[403] = 256'h81FE82990F320837ACDDD50407B888E62518D53E897DACAC5D28BCE8FF3D9339;
        precomp_y[404] = 256'h00E50B1E007B5693C4ECC160D928CD6ED4C978FC6C2A68AFC03F397D72A60383;
        precomp_y[405] = 256'h7D055B74B0195140BC0E2E93A97F07B3A30401487720DF86D3BD18106DF3CC72;
        precomp_y[406] = 256'h1C54A2D39C34B0DB0DEB61B5B5F46033B1E4C58105113BF3D3F38DE1C97CC7E2;
        precomp_y[407] = 256'hB458D7F1390FA4D7D2473863ABEDC063EF310ADF7CA2F2C882BCAD3E02F1B554;
        precomp_y[408] = 256'h8DAAB84B92157D160CA0F160099877A1EF7EF0721BDB5BC689D16A194EBEDEAF;
        precomp_y[409] = 256'h39FFFCB38F74D4719BE8D1A214C61AD3DF4A91BFD599C3AE3B54B4EC0860A942;
        precomp_y[410] = 256'h5BFA8A78D42B95EF327EB0C3692B3BA95EB506A24E2FCA1E391EC54540A76278;
        precomp_y[411] = 256'h6DCB6276CBE37B91162A243F57AFCD9A8CC2C661652C324A567D5DB722A0D750;
        precomp_y[412] = 256'hD1F880AEC18D0191B74578C16D0418F6C7E59F2D157C0D56E25137ECC1B7F74A;
        precomp_y[413] = 256'hF44845811E3266CDF4625390E729154F516947173206EF9B9106C547FF4A21D1;
        precomp_y[414] = 256'hC0550B9A72899A7B42197CFED195C704A6333D5E178D91C10D50B7724140CAD0;
        precomp_y[415] = 256'h1B44E253AF3B214FEDBEB4AC50110DF6D7056D06617C2BF36189A74D64450603;
        precomp_y[416] = 256'h1B5B12A895FB7130E879240674B8F7356730938B675996FBA30A9744960FEBEF;
        precomp_y[417] = 256'h4CC418F82180207EFC846A41ED6973F2814CEB07A8BD252E338E32CDE352EE6F;
        precomp_y[418] = 256'h72946592D3C11404881B972CEBA81D4FF3F80DCD40B15DA5F56E0723841E4F99;
        precomp_y[419] = 256'h5D4AC85189350A54AF58DEF46F3F3D692EF0F6A39DD4EF866BB1101BDF5E6144;
        precomp_y[420] = 256'h56E32E5B8FC2DB2F21D64BAD35E3F11565928533A829D744939BA456BB1774FE;
        precomp_y[421] = 256'h43E4188AC92606C1CD6BEC5BA4EDB0456569F87A625DB932D0F8E71E516B8127;
        precomp_y[422] = 256'h89A7B2C9E9F3588D990F6FA196E366B6054F9A301218A2A9C9B87C4855F0B360;
        precomp_y[423] = 256'h3F03ED1FBE1A661EF43EF9F7D753EAADE3E1A3912A682AD4FB19526CC0011728;
        precomp_y[424] = 256'h38AF8B6130701881FBBFE7245396ADC932C25B84DFBC4DBDA54BD236C04B4FDE;
        precomp_y[425] = 256'h7380D6865F5FD782B0708B3B62C39E49864B2BA74066167CBBCEDE2AB0F84787;
        precomp_y[426] = 256'h4468BF1BEE43F1007E800B68B7B3B2432F3445C5C8ACA59F7534BEAEBB771F41;
        precomp_y[427] = 256'h62777495AE16314FD7D0CEF824A27A9F748C5C9B09C516459C1EC9DD9D7B59F5;
        precomp_y[428] = 256'h2A4EA7DAC87522CB7D92C4508E86D0B939FAD0249FC2CF151BA005CDB743D0BC;
        precomp_y[429] = 256'h07321690DE24499CF52F484089C4D7B411158D52D32731C9FAAEA5678BF6072B;
        precomp_y[430] = 256'h56727C07247B12D6C1ADE4733C69170030E5582ACDE140343449F24159FFA44D;
        precomp_y[431] = 256'h0984DD72855CDEAE7C580046B32CFA7A45B61B75944735E1D5FD9065268AC521;
        precomp_y[432] = 256'hD1593BF5B9E793F725CEA3682CEABB11F06B36AB899E160A0F1F736A80BC9B92;
        precomp_y[433] = 256'h4A89307D27D7F3607ACD1643719BE1481C7EED5C775988838BF6CC13A4723D9F;
        precomp_y[434] = 256'hB5AB61E396F8837628F3389E9999EF55B73A58C0D33DEBC7258125302B96C772;
        precomp_y[435] = 256'h23CCAFAECC84EA723C434342B839CD0AB42173BC1AA1DB201073FE266593403D;
        precomp_y[436] = 256'h03A57F08FFECCCFCCD9A0E7C827D98A2FFCEEA9A6C39D2005CFAE62334EEBA8F;
        precomp_y[437] = 256'hE31161A568D81328C7F9783FDE146D07B51AAE150BFE719D00AB4E9EAE65D172;
        precomp_y[438] = 256'hFAED7EF882733020888EB5305C6DEA4BCACD208F0FBB66B706F3CF41A8864080;
        precomp_y[439] = 256'h287AB9C962126FB7E0340F299EDEB89E7BF235B3B3F08213D630C9DF198ADA1D;
        precomp_y[440] = 256'h95CE721C39929D76B0EA83B180BF25C2E301413D60FB87172E0EE8F0593F8423;
        precomp_y[441] = 256'h18439939496D29A158A532BE76B04932A23E3DDDD51A1B07C6C33E6A11E1AFA8;
        precomp_y[442] = 256'h84CBD8C38DCCF0EFDE3946F3BA2EAC253AAAB9768F7F601E7D95BC74004C7F65;
        precomp_y[443] = 256'hC04C7CC44EA1D8B2273B917019B9EFB36E8F422C4863F718582F57A0778273EE;
        precomp_y[444] = 256'h5BD732642F16D4E77BCC485572494523C221FA1D321C552A53241DD794C7D98E;
        precomp_y[445] = 256'h84439E001571E1EA53BCC24BA11B6F7CDED0A649B2A12FC9C2A618FECB39ADA7;
        precomp_y[446] = 256'hE53840E301110DB189EC241AE7B2CB8929669DA95C07F3D06277F667B90CAD12;
        precomp_y[447] = 256'h9C10F0DBBB16D8074680133FE62E0EAB130CB0B95193785204AFCF4C38814061;
        precomp_y[448] = 256'h3376B6C893AD5EC5991F7EF96A6B11052F2262C6680045FDFC4D4BFEEA64AE75;
        precomp_y[449] = 256'h5E48FCB33ED9C0EC3594EEB0081ADAAABD5EC5A57EEAF01FC9F00D02C692CB06;
        precomp_y[450] = 256'h64496D5085435DE6991A838ED984BC092554053B54B05A2E0490D2CEDA7D5B76;
        precomp_y[451] = 256'h2E1209FBA7921C290E351E6173C02CB5C629D88F04CA51AF30F3712375355213;
        precomp_y[452] = 256'hB2A2CD8B73F76F3D1079198D34441008278F73C893979ECEEEFC59117BA17814;
        precomp_y[453] = 256'h589FC4269466B1FFB9C0CBD4B022E9EE7EDAAE878F4CC240B60DB60D6C28F04F;
        precomp_y[454] = 256'h2D9C53F10EE63B932ADF679D96B548D8D47D8F7458EF8B459664DA23BE32C363;
        precomp_y[455] = 256'hC76852F507159524541569F63C4C9C7D424285E7E83145D5E5161998EFEBF968;
        precomp_y[456] = 256'h88F919BEB9993A1661F78145F54149F46ABFA8591907736DD5E85F25BF2DC7CB;
        precomp_y[457] = 256'h346C98E32BC2A4E8C7689E54EEB1064C1B5691FBCF5A471055CEFBCF18A32F65;
        precomp_y[458] = 256'hD959BDF058D21CC3430527E8CC49DC562DD20BF130F0E13A55CC69CC1E116F35;
        precomp_y[459] = 256'h24F09BBF7BCF50AA0CA239BEB925505E7E99D0FF5A9595745370EEA17B4841F6;
        precomp_y[460] = 256'h9652B4589D269AD968EE7012AEE4744725BA917DF120BDA69D2194EEA56D7B60;
        precomp_y[461] = 256'h8061BB940D6485FED9FBD55766DB3DCAC648C7C42E025494E6C3A91CFD5C609E;
        precomp_y[462] = 256'hAB0C7E38C85EE1CC027964B2DE42372FFD86ECB8FD3F0A8184F5AF3858A7E4EA;
        precomp_y[463] = 256'h08D5B83D0DC3022C04F79723C6F16722CC7EEEB9C964496FC9F67C29351A0BED;
        precomp_y[464] = 256'h0F5868F2C2E872492137339740415C4AECB1F30DB204FE4180E01D79EB536800;
        precomp_y[465] = 256'h5CF10D7403085DD7CC6951453F9F763D6596ABFAEB7CF21634EE07F8A4F141AC;
        precomp_y[466] = 256'h005A90903766D6EBC58C5D609B6A5675E5EC7B7386A17C412574D179A0FD5450;
        precomp_y[467] = 256'h88CF0055ADF1E122535611D7BD3E00A730C9EDD5898D25BFF0ABB9BF6BD6C8C0;
        precomp_y[468] = 256'hC926B3DD0519241D02E776EA16112E41259CE896472CE71FDE4261BD29C678EE;
        precomp_y[469] = 256'hD5B1AADF84D387B8FDDC7B26A7F736A67E296FED7978E81F6E7B3B090E94D733;
        precomp_y[470] = 256'h5358DAF260FEA2A1B9A4C6F1B8BEBE094983499CFE5577A2ED8F817F46B41CCF;
        precomp_y[471] = 256'hDA3C66AFE4CFB3DFF55F67615C6AC42A8DC172415AD38619DFE2A13B7E42FF9E;
        precomp_y[472] = 256'h1098FA7613DCE1C5029F7FEA30740377691AA3CF3D13CF946F2D81912D3B9E83;
        precomp_y[473] = 256'h72724B4D0EEC94DA7494B4D983A2DF06DF96EE83E578D920C25970897B4B3D8A;
        precomp_y[474] = 256'hCDCD21DFE5ED81511A2D8C77E08B76F74939D39F1F5581B0AA9560660FA14A7C;
        precomp_y[475] = 256'hFCD1B2AC39C262C694EEF5E052338F9CCAC2D04DED17C290768759CD13B7D550;
        precomp_y[476] = 256'h143C7DDE0D33BA5BC2AC8D83CC462F942607BFF2A1AA32D9F32E14C282232226;
        precomp_y[477] = 256'h27C341AE87E7AFEEF8AF4598E8E27CABC127B0541B389CFB266EC9D2FE400284;
        precomp_y[478] = 256'hEB642FBBFE3274E52FD1CAE9744FABFAC0DB80E62BD4F7C3FC2CA43B18CE52EF;
        precomp_y[479] = 256'hF5B386DFAC71EB35499D5B2A960FD20E0FDE39FC10DD5C63DC50B55BCD660D9C;
        precomp_y[480] = 256'h504532ED34F97EB9B8B27664AB4400322B8B47F69C403BBD6BC7433016923DEC;
        precomp_y[481] = 256'hA367B5844F9B7B2BA82FCCCAB9A12A8C2C1CA5F73E630173E37E600F0F2FCFB6;
        precomp_y[482] = 256'h90B0CD33C350EA2E54C252647A3FC91F5B4F9DC31F58E86FC47825DCE3D0F43A;
        precomp_y[483] = 256'h17E38880F10B9927764C4997326B0B9F63D0E03A0FD2F0BDB1FF3CCA1F566BB7;
        precomp_y[484] = 256'h66BB180A7EAA64D84BFE6A17D457F5E7073964ACFF9087293BC540AA1CB6464F;
        precomp_y[485] = 256'hE208BE8A88BE7B3F6B6B06CEA3AAFB45C439F0BAD517A784BA13F80B707CAF14;
        precomp_y[486] = 256'hF8029F31B8E5EE3F77A758AE343BE25834C7BEF4C1B555C74CB63D51CBA5FEC1;
        precomp_y[487] = 256'hE4ABD7F9FE40F27D5B7B76516A9FD714AACD2AE05F0A1F10E94327E376F0AF52;
        precomp_y[488] = 256'h81E9997A8B1C594906554BCF154166D340F9EA5FCE55EC83EED793D55CA3E513;
        precomp_y[489] = 256'h7837965ECF26A7F3428D286441E1D09A91EAFF0C5ECD2C28BC81776667FA35B1;
        precomp_y[490] = 256'h72688262594C75BBBB55C0FAAF7991C8F412E0EB0AFD1C0CF5BCAB82D8DAF31A;
        precomp_y[491] = 256'h479FC222A7BCAA62AEE807C4BA6309E6CFBCC783AFD49ECC0FB9B45FCF84673D;
        precomp_y[492] = 256'h1C965FE7A82190529D25EE0CE1FD62F37196431D7BD78302E287A26A2EEAA23E;
        precomp_y[493] = 256'hBB79E77224B02FCFDD1E3C9CEDBAD212EA875C751FE7C81E76D7D0D9A372236E;
        precomp_y[494] = 256'hD0D978424F0010A40DF9EB8B8E5D8147F618DA4374B8A4DB222E4AB2B32B3D92;
        precomp_y[495] = 256'h60B66D45A693175A3A38BB4FEFB32DAC1CB558E1B0D13571E24A14D59452BDC0;
        precomp_y[496] = 256'hEB3BD91E9C09178A398E112A9264484EC1980C19B1993B13560D39FB92295F7A;
        precomp_y[497] = 256'hBB507868C1E0528251B635B9DCF28E5AC5770C05C7AFC2A3F4B4C45B7D8993EC;
        precomp_y[498] = 256'hCC99452B85092CA539CC1B6683B7AB371B8A6525269A1ECF91B857BEE1DB3BD4;
        precomp_y[499] = 256'hDDAC2D377F03C201FFA0419D6596D10327D6C70313BB492FF495F946285D8F38;
        precomp_y[500] = 256'hF21EE70050DBB61C238C89E62942353871B010E798867BDD149AD28B3F28CADF;
        precomp_y[501] = 256'h8BC13ECC207EFD91F7F4C4426E9A425AA17B557820404ECAB09D5582D41F7379;
        precomp_y[502] = 256'h5DC23258F93D7DB5E5799195B74E95194C300A9128F924C1C1E4865E02D8407D;
        precomp_y[503] = 256'h720A8104473DC90465585ED21A0244F0FBB5A2865B8E51175A21F6448776BB7B;
        precomp_y[504] = 256'hF729D335210E80618A8ABDCDB71AABE193F50ADADFAF7D52783991DDD3CA5D4B;
        precomp_y[505] = 256'h9649994D64705B8762C98BBF1B41B7252B814A893E780FDF5689C9DA0692D6FF;
        precomp_y[506] = 256'h868B3E4F9AE4BEA8EFDE50BFC5A5B2680B74B4A874E86DE6E9AE476F10B3B778;
        precomp_y[507] = 256'h01ABA673D0372029546C174A3A72268CEE9D7E41DD97DE2FFCBE1F9F1A5288B9;
        precomp_y[508] = 256'hD90E94ECB50BFEE8C951AFB8E65C7386875EA99E31F553E866E0034206D39698;
        precomp_y[509] = 256'hEBFE58495A1E6A3646C382208656F638ED0AEC0AD40C0524017071023126F795;
        precomp_y[510] = 256'hD36AE886A0ACBC9AD1564D974D3F0309E9039B93BB350D922B7F8C7AC6BFA042;
        precomp_y[511] = 256'h1298FDD70E448D2D799863026B4B2D4902B32148D6D1E5F815F5B0C005C9E21F;
    end

    // -----------------------------
    // Operações de curva (já existentes no seu projeto)
    // -----------------------------
    reg         dbl_start;
    wire [255:0] dbl_x, dbl_y, dbl_z;
    wire        dbl_done;

    reg         add_start;
    reg [255:0] add_px, add_py;
    wire [255:0] add_x, add_y, add_z;
    wire        add_done;

    reg         inv_start;
    wire [255:0] inv_out;
    wire        inv_done;

    reg         mul_start;
    reg [255:0] mul_a, mul_b;
    wire [255:0] mul_result;
    wire        mul_done;
    reg [255:0] rx, ry, rz;
    secp256k1_point_double u_double (
        .clk(clk), .rst_n(rst_n), .start(dbl_start),
        .x1(rx), .y1(ry), .z1(rz),
        .x3(dbl_x), .y3(dbl_y), .z3(dbl_z),
        .done(dbl_done)
    );

    secp256k1_point_add u_add (
        .clk(clk), .rst_n(rst_n), .start(add_start),
        .x1(rx), .y1(ry), .z1(rz),
        .x2(add_px), .y2(add_py),
        .x3(add_x), .y3(add_y), .z3(add_z),
        .done(add_done)
    );

    secp256k1_inv_mod u_inv (
        .clk(clk), .rst_n(rst_n), .start(inv_start),
        .a(rz), .result(inv_out), .done(inv_done)
    );

    secp256k1_mul_mod u_mul (
        .clk(clk), .rst_n(rst_n), .start(mul_start),
        .a(mul_a), .b(mul_b), .result(mul_result), .done(mul_done)
    );

    // -----------------------------
    // Acumulador Jacobiano
    // -----------------------------

    reg         r_is_inf;

    // -----------------------------
    // wNAF storage (RAM de bytes)
    // -----------------------------
    localparam integer NAF_LEN = 264;
	reg  [7:0] naf_mem [0:NAF_LEN-1];



    reg [264:0] naf_k;
    reg [8:0]   naf_bit_pos;
    reg [8:0]   naf_len;
    reg [8:0]   digit_pos;

    // leitura síncrona do byte atual (evita mux gigante)
    reg [8:0]         naf_addr;
    reg signed [7:0]  naf_q;
    always @(posedge clk) begin
        naf_q <= naf_mem[naf_addr];
    end

    reg found_first;

    // Flags de espera
    reg wait_dbl, wait_add, wait_inv, wait_mul;

    // Afim
    reg [255:0] z_inv, z2, z3;

    // -----------------------------
    // FSM
    // -----------------------------
    reg [4:0] state;

    localparam IDLE        = 5'd0;
    localparam INIT        = 5'd1;
    localparam CONVERT_NAF = 5'd2;
    localparam WAIT_NAF    = 5'd3;
    localparam FIND_MSB    = 5'd4;
    localparam DOUBLE      = 5'd5;
    localparam WAIT_DOUBLE = 5'd6;
    localparam CHECK_DIGIT = 5'd7;
    localparam WAIT_ROM    = 5'd8;
    localparam ADD_POINT   = 5'd9;
    localparam WAIT_ADD    = 5'd10;
    localparam NEXT_DIGIT  = 5'd11;
    localparam TO_AFFINE   = 5'd12;
    localparam WAIT_INV    = 5'd13;
    localparam CALC_Z2     = 5'd14;
    localparam CALC_QX     = 5'd15;
    localparam CALC_Z3     = 5'd16;
    localparam CALC_QY     = 5'd17;
    localparam DONE_STATE  = 5'd18;

    // -----------------------------
    // FSM sequencial
    // -----------------------------
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            qx <= 256'd0; qy <= 256'd0;
            done <= 1'b0;
            point_at_inf <= 1'b0;

            rx <= 256'd0; ry <= 256'd0; rz <= 256'd0;
            r_is_inf <= 1'b1;

            state <= IDLE;

            naf_k <= 265'd0;
            naf_bit_pos <= 9'd0;
            naf_len <= 9'd0;
            digit_pos <= 9'd0;
            naf_addr <= 9'd0;
            naf_q <= 8'sd0;

            found_first <= 1'b0;

            dbl_start <= 1'b0;
            add_start <= 1'b0;
            inv_start <= 1'b0;
            mul_start <= 1'b0;

            wait_dbl <= 1'b0;
            wait_add <= 1'b0;
            wait_inv <= 1'b0;
            wait_mul <= 1'b0;

            rom_addr <= 'b0;
            rom_neg <= 1'b0;
            rom_wait <= 1'b0;
            rom_use_add <= 1'b0;

            add_px <= 256'd0;
            add_py <= 256'd0;

            z_inv <= 256'd0;
            z2 <= 256'd0;
            z3 <= 256'd0;

        end else begin
            // defaults
            done      <= 1'b0;
            dbl_start <= 1'b0;
            add_start <= 1'b0;
            inv_start <= 1'b0;
            mul_start <= 1'b0;

            case (state)
                IDLE: begin
                    point_at_inf <= 1'b0;
                    if (start) begin
                        // este core "barato" assume use_g=1 (tabela fixa)
                        if (!use_g) begin
                            $display("AVISO: use_g=0 ignorado neste core (tabela fixa do G).");
                        end

                        if (k == 256'd0) begin
                            point_at_inf <= 1'b1;
                            qx <= 256'd0;
                            qy <= 256'd0;
                            state <= DONE_STATE;
                        end else begin
                            state <= INIT;
                        end
                    end
                end

                INIT: begin
                    naf_k       <= {9'd0, k};
                    naf_bit_pos <= 9'd0;
                    naf_len     <= 9'd0;

                    rx <= 256'd0; ry <= 256'd0; rz <= 256'd0;
                    r_is_inf <= 1'b1;
                    found_first <= 1'b0;

                    state <= CONVERT_NAF;
                end

                CONVERT_NAF: begin : CONV_BLK
                    // constantes
                    reg [264:0] pow2w_ext;
                    reg [W-1:0] wnd;
                    reg [W-1:0] halfw;
                    reg signed [8:0] digit_s;
                    reg [264:0] k_adj;

                    pow2w_ext = (265'd1 << W);
                    halfw = (1 << (W-1));

                    if (naf_k == 265'd0) begin
                        naf_len <= naf_bit_pos;
                        state   <= FIND_MSB;

                    end else if (naf_bit_pos >= NAF_LEN) begin
                        naf_len <= NAF_LEN;
                        state   <= FIND_MSB;

                    end else if (naf_k[0]) begin
                        wnd = naf_k[W-1:0];

                        if (wnd >= halfw) begin
                            digit_s = $signed({1'b0, wnd}) - $signed(pow2w_ext[8:0]); // negativo
                            naf_mem[naf_bit_pos] <= digit_s[7:0];
                            k_adj = naf_k + (pow2w_ext - {{(265-W){1'b0}}, wnd});
                        end else begin
                            digit_s = $signed({1'b0, wnd});
                            naf_mem[naf_bit_pos] <= digit_s[7:0];
                            k_adj = naf_k - {{(265-W){1'b0}}, wnd};
                        end

                        naf_k       <= (k_adj >> 1);
                        naf_bit_pos <= naf_bit_pos + 1'b1;

                    end else begin
                        naf_mem[naf_bit_pos] <= 8'sd0;
                        naf_k       <= (naf_k >> 1);
                        naf_bit_pos <= naf_bit_pos + 1'b1;
                    end
                end

                FIND_MSB: begin
                    if (naf_len == 9'd0) begin
                        point_at_inf <= 1'b1;
                        qx <= 256'd0;
                        qy <= 256'd0;
                        state <= DONE_STATE;
                    end else begin
                        digit_pos <= naf_len - 1'b1;
                        naf_addr  <= naf_len - 1'b1; // 1 ciclo pra ler
                        r_is_inf <= 1'b1;
                        found_first <= 1'b0;
                        state <= WAIT_NAF;
                    end
                end

                WAIT_NAF: begin
                    state <= CHECK_DIGIT;
                end

                DOUBLE: begin
                    // já deixamos o naf_addr apontando pro próximo dígito no NEXT_DIGIT
                    if (!r_is_inf) begin
                        dbl_start <= 1'b1;
                        wait_dbl  <= 1'b1;
                        state     <= WAIT_DOUBLE;
                    end else begin
                        state <= CHECK_DIGIT;
                    end
                end

                WAIT_DOUBLE: begin
                    if (wait_dbl && dbl_done) begin
                        wait_dbl <= 1'b0;
                        rx <= dbl_x;
                        ry <= dbl_y;
                        rz <= dbl_z;
                        state <= CHECK_DIGIT;
                    end
                end

                CHECK_DIGIT: begin : CD_BLK
                    reg signed [8:0] d;
                    reg [8:0]        ad;

                    d  = naf_q;
                    if (d == 0) begin
                        state <= NEXT_DIGIT;
                    end else begin
                        ad = (d < 0) ? -d : d;

                        // idx = (|d|-1)/2  => 0..(NUM_POINTS-1)
                        rom_addr    <= (ad - 1) >> 1;
                        rom_neg     <= (d < 0);
                        rom_use_add <= found_first; // se já iniciou => ADD, senão INIT
                        rom_wait    <= 1'b1;
                        state       <= WAIT_ROM;
                    end
                end

                WAIT_ROM: begin
                    if (rom_wait) begin
                        rom_wait <= 1'b0;
                    end else begin
                        if (!rom_use_add) begin
                            // INIT acumulador
                            rx <= rom_x_q;
                            ry <= rom_neg ? (SECP256K1_P - rom_y_q) : rom_y_q;
                            rz <= 256'd1;
                            r_is_inf <= 1'b0;
                            found_first <= 1'b1;
                            state <= NEXT_DIGIT;
                        end else begin
                            // preparar add
                            add_px <= rom_x_q;
                            add_py <= rom_neg ? (SECP256K1_P - rom_y_q) : rom_y_q;
                            state  <= ADD_POINT;
                        end
                    end
                end

                ADD_POINT: begin
                    if (r_is_inf) begin
                        rx <= add_px;
                        ry <= add_py;
                        rz <= 256'd1;
                        r_is_inf <= 1'b0;
                        state <= NEXT_DIGIT;
                    end else begin
                        add_start <= 1'b1;
                        wait_add  <= 1'b1;
                        state     <= WAIT_ADD;
                    end
                end

                WAIT_ADD: begin
                    if (wait_add && add_done) begin
                        wait_add <= 1'b0;
                        rx <= add_x;
                        ry <= add_y;
                        rz <= add_z;
                        state <= NEXT_DIGIT;
                    end
                end

                NEXT_DIGIT: begin
                    if (digit_pos == 9'd0) begin
                        if (r_is_inf) begin
                            point_at_inf <= 1'b1;
                            qx <= 256'd0;
                            qy <= 256'd0;
                            state <= DONE_STATE;
                        end else begin
                            state <= TO_AFFINE;
                        end
                    end else begin
                        digit_pos <= digit_pos - 1'b1;
                        naf_addr  <= digit_pos - 1'b1; // prefetch do próximo dígito
                        state <= DOUBLE;
                    end
                end

                TO_AFFINE: begin
                    if (rz == 256'd0) begin
                        point_at_inf <= 1'b1;
                        qx <= 256'd0;
                        qy <= 256'd0;
                        state <= DONE_STATE;
                    end else begin
                        inv_start <= 1'b1;
                        wait_inv  <= 1'b1;
                        state     <= WAIT_INV;
                    end
                end

                WAIT_INV: begin
                    if (wait_inv && inv_done) begin
                        wait_inv <= 1'b0;
                        z_inv <= inv_out;

                        mul_a <= inv_out;
                        mul_b <= inv_out;
                        mul_start <= 1'b1;
                        wait_mul  <= 1'b1;
                        state <= CALC_Z2;
                    end
                end

                CALC_Z2: begin
                    if (wait_mul && mul_done) begin
                        wait_mul <= 1'b0;
                        z2 <= mul_result;

                        mul_a <= rx;
                        mul_b <= mul_result;
                        mul_start <= 1'b1;
                        wait_mul  <= 1'b1;
                        state <= CALC_QX;
                    end
                end

                CALC_QX: begin
                    if (wait_mul && mul_done) begin
                        wait_mul <= 1'b0;
                        qx <= mul_result;

                        mul_a <= z2;
                        mul_b <= z_inv;
                        mul_start <= 1'b1;
                        wait_mul  <= 1'b1;
                        state <= CALC_Z3;
                    end
                end

                CALC_Z3: begin
                    if (wait_mul && mul_done) begin
                        wait_mul <= 1'b0;
                        z3 <= mul_result;

                        mul_a <= ry;
                        mul_b <= mul_result;
                        mul_start <= 1'b1;
                        wait_mul  <= 1'b1;
                        state <= CALC_QY;
                    end
                end

                CALC_QY: begin
                    if (wait_mul && mul_done) begin
                        wait_mul <= 1'b0;
                        qy <= mul_result;
                        state <= DONE_STATE;
                    end
                end

                DONE_STATE: begin
                    done  <= 1'b1;
                    state <= IDLE;
                end

                default: state <= IDLE;
            endcase
        end
    end

endmodule
