precomp_x[0] = 256'h79BE667EF9DCBBAC55A06295CE870B07029BFCDB2DCE28D959F2815B16F81798;
precomp_x[1] = 256'hF9308A019258C31049344F85F89D5229B531C845836F99B08601F113BCE036F9;
precomp_x[2] = 256'h2F8BDE4D1A07209355B4A7250A5C5128E88B84BDDC619AB7CBA8D569B240EFE4;
precomp_x[3] = 256'h5CBDF0646E5DB4EAA398F365F2EA7A0E3D419B7E0330E39CE92BDDEDCAC4F9BC;
precomp_x[4] = 256'hACD484E2F0C7F65309AD178A9F559ABDE09796974C57E714C35F110DFC27CCBE;
precomp_x[5] = 256'h774AE7F858A9411E5EF4246B70C65AAC5649980BE5C17891BBEC17895DA008CB;
precomp_x[6] = 256'hF28773C2D975288BC7D1D205C3748651B075FBC6610E58CDDEEDDF8F19405AA8;
precomp_x[7] = 256'hD7924D4F7D43EA965A465AE3095FF41131E5946F3C85F79E44ADBCF8E27E080E;
precomp_x[8] = 256'hDEFDEA4CDB677750A420FEE807EACF21EB9898AE79B9768766E4FAA04A2D4A34;
precomp_x[9] = 256'h2B4EA0A797A443D293EF5CFF444F4979F06ACFEBD7E86D277475656138385B6C;
precomp_x[10] = 256'h352BBF4A4CDD12564F93FA332CE333301D9AD40271F8107181340AEF25BE59D5;
precomp_x[11] = 256'h2FA2104D6B38D11B0230010559879124E42AB8DFEFF5FF29DC9CDADD4ECACC3F;
precomp_x[12] = 256'h9248279B09B4D68DAB21A9B066EDDA83263C3D84E09572E269CA0CD7F5453714;
precomp_x[13] = 256'hDAED4F2BE3A8BF278E70132FB0BEB7522F570E144BF615C07E996D443DEE8729;
precomp_x[14] = 256'hC44D12C7065D812E8ACF28D7CBB19F9011ECD9E9FDF281B0E6A3B5E87D22E7DB;
precomp_x[15] = 256'h6A245BF6DC698504C89A20CFDED60853152B695336C28063B61C65CBD269E6B4;
precomp_x[16] = 256'h1697FFA6FD9DE627C077E3D2FE541084CE13300B0BEC1146F95AE57F0D0BD6A5;
precomp_x[17] = 256'h605BDB019981718B986D0F07E834CB0D9DEB8360FFB7F61DF982345EF27A7479;
precomp_x[18] = 256'h62D14DAB4150BF497402FDC45A215E10DCB01C354959B10CFE31C7E9D87FF33D;
precomp_x[19] = 256'h80C60AD0040F27DADE5B4B06C408E56B2C50E9F56B9B8B425E555C2F86308B6F;
precomp_x[20] = 256'h7A9375AD6167AD54AA74C6348CC54D344CC5DC9487D847049D5EABB0FA03C8FB;
precomp_x[21] = 256'hD528ECD9B696B54C907A9ED045447A79BB408EC39B68DF504BB51F459BC3FFC9;
precomp_x[22] = 256'h049370A4B5F43412EA25F514E8ECDAD05266115E4A7ECB1387231808F8B45963;
precomp_x[23] = 256'h77F230936EE88CBBD73DF930D64702EF881D811E0E1498E2F1C13EB1FC345D74;
precomp_x[24] = 256'hF2DAC991CC4CE4B9EA44887E5C7C0BCE58C80074AB9D4DBAEB28531B7739F530;
precomp_x[25] = 256'h463B3D9F662621FB1B4BE8FBBE2520125A216CDFC9DAE3DEBCBA4850C690D45B;
precomp_x[26] = 256'hF16F804244E46E2A09232D4AFF3B59976B98FAC14328A2D1A32496B49998F247;
precomp_x[27] = 256'hCAF754272DC84563B0352B7A14311AF55D245315ACE27C65369E15F7151D41D1;
precomp_x[28] = 256'h2600CA4B282CB986F85D0F1709979D8B44A09C07CB86D7C124497BC86F082120;
precomp_x[29] = 256'h7635CA72D7E8432C338EC53CD12220BC01C48685E24F7DC8C602A7746998E435;
precomp_x[30] = 256'h754E3239F325570CDBBF4A87DEEE8A66B7F2B33479D468FBC1A50743BF56CC18;
precomp_x[31] = 256'hE3E6BD1071A1E96AFF57859C82D570F0330800661D1C952F9FE2694691D9B9E8;
precomp_x[32] = 256'h186B483D056A033826AE73D88F732985C4CCB1F32BA35F4B4CC47FDCF04AA6EB;
precomp_x[33] = 256'hDF9D70A6B9876CE544C98561F4BE4F725442E6D2B737D9C91A8321724CE0963F;
precomp_x[34] = 256'h5EDD5CC23C51E87A497CA815D5DCE0F8AB52554F849ED8995DE64C5F34CE7143;
precomp_x[35] = 256'h290798C2B6476830DA12FE02287E9E777AA3FBA1C355B17A722D362F84614FBA;
precomp_x[36] = 256'hAF3C423A95D9F5B3054754EFA150AC39CD29552FE360257362DFDECEF4053B45;
precomp_x[37] = 256'h766DBB24D134E745CCCAA28C99BF274906BB66B26DCF98DF8D2FED50D884249A;
precomp_x[38] = 256'h59DBF46F8C94759BA21277C33784F41645F7B44F6C596A58CE92E666191ABE3E;
precomp_x[39] = 256'hF13ADA95103C4537305E691E74E9A4A8DD647E711A95E73CB62DC6018CFD87B8;
precomp_x[40] = 256'h7754B4FA0E8ACED06D4167A2C59CCA4CDA1869C06EBADFB6488550015A88522C;
precomp_x[41] = 256'h948DCADF5990E048AA3874D46ABEF9D701858F95DE8041D2A6828C99E2262519;
precomp_x[42] = 256'h7962414450C76C1689C7B48F8202EC37FB224CF5AC0BFA1570328A8A3D7C77AB;
precomp_x[43] = 256'h3514087834964B54B15B160644D915485A16977225B8847BB0DD085137EC47CA;
precomp_x[44] = 256'hD3CC30AD6B483E4BC79CE2C9DD8BC54993E947EB8DF787B442943D3F7B527EAF;
precomp_x[45] = 256'h1624D84780732860CE1C78FCBFEFE08B2B29823DB913F6493975BA0FF4847610;
precomp_x[46] = 256'h733CE80DA955A8A26902C95633E62A985192474B5AF207DA6DF7B4FD5FC61CD4;
precomp_x[47] = 256'h15D9441254945064CF1A1C33BBD3B49F8966C5092171E699EF258DFAB81C045C;
precomp_x[48] = 256'hA1D0FCF2EC9DE675B612136E5CE70D271C21417C9D2B8AAAAC138599D0717940;
precomp_x[49] = 256'hE22FBE15C0AF8CCC5780C0735F84DBE9A790BADEE8245C06C7CA37331CB36980;
precomp_x[50] = 256'h311091DD9860E8E20EE13473C1155F5F69635E394704EAA74009452246CFA9B3;
precomp_x[51] = 256'h34C1FD04D301BE89B31C0442D3E6AC24883928B45A9340781867D4232EC2DBDF;
precomp_x[52] = 256'hF219EA5D6B54701C1C14DE5B557EB42A8D13F3ABBCD08AFFCC2A5E6B049B8D63;
precomp_x[53] = 256'hD7B8740F74A8FBAAB1F683DB8F45DE26543A5490BCA627087236912469A0B448;
precomp_x[54] = 256'h32D31C222F8F6F0EF86F7C98D3A3335EAD5BCD32ABDD94289FE4D3091AA824BF;
precomp_x[55] = 256'h7461F371914AB32671045A155D9831EA8793D77CD59592C4340F86CBC18347B5;
precomp_x[56] = 256'hEE079ADB1DF1860074356A25AA38206A6D716B2C3E67453D287698BAD7B2B2D6;
precomp_x[57] = 256'h16EC93E447EC83F0467B18302EE620F7E65DE331874C9DC72BFD8616BA9DA6B5;
precomp_x[58] = 256'hEAA5F980C245F6F038978290AFA70B6BD8855897F98B6AA485B96065D537BD99;
precomp_x[59] = 256'h078C9407544AC132692EE1910A02439958AE04877151342EA96C4B6B35A49F51;
precomp_x[60] = 256'h494F4BE219A1A77016DCD838431AEA0001CDC8AE7A6FC688726578D9702857A5;
precomp_x[61] = 256'hA598A8030DA6D86C6BC7F2F5144EA549D28211EA58FAA70EBF4C1E665C1FE9B5;
precomp_x[62] = 256'hC41916365ABB2B5D09192F5F2DBEAFEC208F020F12570A184DBADC3E58595997;
precomp_x[63] = 256'h841D6063A586FA475A724604DA03BC5B92A2E0D2E0A36ACFE4C73A5514742881;
precomp_x[64] = 256'h5E95BB399A6971D376026947F89BDE2F282B33810928BE4DED112AC4D70E20D5;
precomp_x[65] = 256'h36E4641A53948FD476C39F8A99FD974E5EC07564B5315D8BF99471BCA0EF2F66;
precomp_x[66] = 256'h0336581EA7BFBBB290C191A2F507A41CF5643842170E914FAEAB27C2C579F726;
precomp_x[67] = 256'h8AB89816DADFD6B6A1F2634FCF00EC8403781025ED6890C4849742706BD43EDE;
precomp_x[68] = 256'h1E33F1A746C9C5778133344D9299FCAA20B0938E8ACFF2544BB40284B8C5FB94;
precomp_x[69] = 256'h85B7C1DCB3CEC1B7EE7F30DED79DD20A0ED1F4CC18CBCFCFA410361FD8F08F31;
precomp_x[70] = 256'h29DF9FBD8D9E46509275F4B125D6D45D7FBE9A3B878A7AF872A2800661AC5F51;
precomp_x[71] = 256'hA0B1CAE06B0A847A3FEA6E671AAF8ADFDFE58CA2F768105C8082B2E449FCE252;
precomp_x[72] = 256'h04E8CEAFB9B3E9A136DC7FF67E840295B499DFB3B2133E4BA113F2E4C0E121E5;
precomp_x[73] = 256'hD24A44E047E19B6F5AFB81C7CA2F69080A5076689A010919F42725C2B789A33B;
precomp_x[74] = 256'hEA01606A7A6C9CDD249FDFCFACB99584001EDD28ABBAB77B5104E98E8E3B35D4;
precomp_x[75] = 256'hAF8ADDBF2B661C8A6C6328655EB96651252007D8C5EA31BE4AD196DE8CE2131F;
precomp_x[76] = 256'h00E3AE1974566CA06CC516D47E0FB165A674A3DABCFCA15E722F0E3450F45889;
precomp_x[77] = 256'h591EE355313D99721CF6993FFED1E3E301993FF3ED258802075EA8CED397E246;
precomp_x[78] = 256'h11396D55FDA54C49F19AA97318D8DA61FA8584E47B084945077CF03255B52984;
precomp_x[79] = 256'h3C5D2A1BA39C5A1790000738C9E0C40B8DCDFD5468754B6405540157E017AA7A;
precomp_x[80] = 256'hCC8704B8A60A0DEFA3A99A7299F2E9C3FBC395AFB04AC078425EF8A1793CC030;
precomp_x[81] = 256'hC533E4F7EA8555AACD9777AC5CAD29B97DD4DEFCCC53EE7EA204119B2889B197;
precomp_x[82] = 256'h0C14F8F2CCB27D6F109F6D08D03CC96A69BA8C34EEC07BBCF566D48E33DA6593;
precomp_x[83] = 256'hA6CBC3046BC6A450BAC24789FA17115A4C9739ED75F8F21CE441F72E0B90E6EF;
precomp_x[84] = 256'h347D6D9A02C48927EBFB86C1359B1CAF130A3C0267D11CE6344B39F99D43CC38;
precomp_x[85] = 256'hDA6545D2181DB8D983F7DCB375EF5866D47C67B1BF31C8CF855EF7437B72656A;
precomp_x[86] = 256'hC40747CC9D012CB1A13B8148309C6DE7EC25D6945D657146B9D5994B8FEB1111;
precomp_x[87] = 256'h4E42C8EC82C99798CCF3A610BE870E78338C7F713348BD34C8203EF4037F3502;
precomp_x[88] = 256'h3775AB7089BC6AF823ABA2E1AF70B236D251CADB0C86743287522A1B3B0DEDEA;
precomp_x[89] = 256'hCEE31CBF7E34EC379D94FB814D3D775AD954595D1314BA8846959E3E82F74E26;
precomp_x[90] = 256'hB4F9EAEA09B6917619F6EA6A4EB5464EFDDB58FD45B1EBEFCDC1A01D08B47986;
precomp_x[91] = 256'hD4263DFC3D2DF923A0179A48966D30CE84E2515AFC3DCCC1B77907792EBCC60E;
precomp_x[92] = 256'h48457524820FA65A4F8D35EB6930857C0032ACC0A4A2DE422233EEDA897612C4;
precomp_x[93] = 256'hDFEEEF1881101F2CB11644F3A2AFDFC2045E19919152923F367A1767C11CCEDA;
precomp_x[94] = 256'h6D7EF6B17543F8373C573F44E1F389835D89BCBC6062CED36C82DF83B8FAE859;
precomp_x[95] = 256'hE75605D59102A5A2684500D3B991F2E3F3C88B93225547035AF25AF66E04541F;
precomp_x[96] = 256'hEB98660F4C4DFAA06A2BE453D5020BC99A0C2E60ABE388457DD43FEFB1ED620C;
precomp_x[97] = 256'h13E87B027D8514D35939F2E6892B19922154596941888336DC3563E3B8DBA942;
precomp_x[98] = 256'hEE163026E9FD6FE017C38F06A5BE6FC125424B371CE2708E7BF4491691E5764A;
precomp_x[99] = 256'hB268F5EF9AD51E4D78DE3A750C2DC89B1E626D43505867999932E5DB33AF3D80;
precomp_x[100] = 256'hFF07F3118A9DF035E9FAD85EB6C7BFE42B02F01CA99CEEA3BF7FFDBA93C4750D;
precomp_x[101] = 256'h8D8B9855C7C052A34146FD20FFB658BEA4B9F69E0D825EBEC16E8C3CE2B526A1;
precomp_x[102] = 256'h52DB0B5384DFBF05BFA9D472D7AE26DFE4B851CECA91B1EBA54263180DA32B63;
precomp_x[103] = 256'hE62F9490D3D51DA6395EFD24E80919CC7D0F29C3F3FA48C6FFF543BECBD43352;
precomp_x[104] = 256'h7F30EA2476B399B4957509C88F77D0191AFA2FF5CB7B14FD6D8E7D65AAAB1193;
precomp_x[105] = 256'h5098FF1E1D9F14FB46A210FADA6C903FEF0FB7B4A1DD1D9AC60A0361800B7A00;
precomp_x[106] = 256'h32B78C7DE9EE512A72895BE6B9CBEFA6E2F3C4CCCE445C96B9F2C81E2778AD58;
precomp_x[107] = 256'hE2CB74FDDC8E9FBCD076EEF2A7C72B0CE37D50F08269DFC074B581550547A4F7;
precomp_x[108] = 256'h8438447566D4D7BEDADC299496AB357426009A35F235CB141BE0D99CD10AE3A8;
precomp_x[109] = 256'h4162D488B89402039B584C6FC6C308870587D9C46F660B878AB65C82C711D67E;
precomp_x[110] = 256'h3FAD3FA84CAF0F34F0F89BFD2DCF54FC175D767AEC3E50684F3BA4A4BF5F683D;
precomp_x[111] = 256'h674F2600A3007A00568C1A7CE05D0816C1FB84BF1370798F1C69532FAEB1A86B;
precomp_x[112] = 256'hD32F4DA54ADE74ABB81B815AD1FB3B263D82D6C692714BCFF87D29BD5EE9F08F;
precomp_x[113] = 256'h30E4E670435385556E593657135845D36FBB6931F72B08CB1ED954F1E3CE3FF6;
precomp_x[114] = 256'hBE2062003C51CC3004682904330E4DEE7F3DCD10B01E580BF1971B04D4CAD297;
precomp_x[115] = 256'h93144423ACE3451ED29E0FB9AC2AF211CB6E84A601DF5993C419859FFF5DF04A;
precomp_x[116] = 256'hB015F8044F5FCBDCF21CA26D6C34FB8197829205C7B7D2A7CB66418C157B112C;
precomp_x[117] = 256'hD5E9E1DA649D97D89E4868117A465A3A4F8A18DE57A140D36B3F2AF341A21B52;
precomp_x[118] = 256'hD3AE41047DD7CA065DBF8ED77B992439983005CD72E16D6F996A5316D36966BB;
precomp_x[119] = 256'h463E2763D885F958FC66CDD22800F0A487197D0A82E377B49F80AF87C897B065;
precomp_x[120] = 256'h7985FDFD127C0567C6F53EC1BB63EC3158E597C40BFE747C83CDDFC910641917;
precomp_x[121] = 256'h74A1AD6B5F76E39DB2DD249410EAC7F99E74C59CB83D2D0ED5FF1543DA7703E9;
precomp_x[122] = 256'h30682A50703375F602D416664BA19B7FC9BAB42C72747463A71D0896B22F6DA3;
precomp_x[123] = 256'h9E2158F0D7C0D5F26C3791EFEFA79597654E7A2B2464F52B1EE6C1347769EF57;
precomp_x[124] = 256'h176E26989A43C9CFEBA4029C202538C28172E566E3C4FCE7322857F3BE327D66;
precomp_x[125] = 256'h75D46EFEA3771E6E68ABB89A13AD747ECF1892393DFC4F1B7004788C50374DA8;
precomp_x[126] = 256'h809A20C67D64900FFB698C4C825F6D5F2310FB0451C869345B7319F645605721;
precomp_x[127] = 256'h1B38903A43F7F114ED4500B4EAC7083FDEFECE1CF29C63528D563446F972C180;
precomp_y[0] = 256'h483ADA7726A3C4655DA4FBFC0E1108A8FD17B448A68554199C47D08FFB10D4B8;
precomp_y[1] = 256'h388F7B0F632DE8140FE337E62A37F3566500A99934C2231B6CB9FD7584B8E672;
precomp_y[2] = 256'hD8AC222636E5E3D6D4DBA9DDA6C9C426F788271BAB0D6840DCA87D3AA6AC62D6;
precomp_y[3] = 256'h6AEBCA40BA255960A3178D6D861A54DBA813D0B813FDE7B5A5082628087264DA;
precomp_y[4] = 256'hCC338921B0A7D9FD64380971763B61E9ADD888A4375F8E0F05CC262AC64F9C37;
precomp_y[5] = 256'hD984A032EB6B5E190243DD56D7B7B365372DB1E2DFF9D6A8301D74C9C953C61B;
precomp_y[6] = 256'h0AB0902E8D880A89758212EB65CDAF473A1A06DA521FA91F29B5CB52DB03ED81;
precomp_y[7] = 256'h581E2872A86C72A683842EC228CC6DEFEA40AF2BD896D3A5C504DC9FF6A26B58;
precomp_y[8] = 256'h4211AB0694635168E997B0EAD2A93DAECED1F4A04A95C0F6CFB199F69E56EB77;
precomp_y[9] = 256'h85E89BC037945D93B343083B5A1C86131A01F60C50269763B570C854E5C09B7A;
precomp_y[10] = 256'h321EB4075348F534D59C18259DDA3E1F4A1B3B2E71B1039C67BD3D8BCF81998C;
precomp_y[11] = 256'h02DE1068295DD865B64569335BD5DD80181D70ECFC882648423BA76B532B7D67;
precomp_y[12] = 256'h73016F7BF234AADE5D1AA71BDEA2B1FF3FC0DE2A887912FFE54A32CE97CB3402;
precomp_y[13] = 256'hA69DCE4A7D6C98E8D4A1ACA87EF8D7003F83C230F3AFA726AB40E52290BE1C55;
precomp_y[14] = 256'h2119A460CE326CDC76C45926C982FDAC0E106E861EDF61C5A039063F0E0E6482;
precomp_y[15] = 256'hE022CF42C2BD4A708B3F5126F16A24AD8B33BA48D0423B6EFD5E6348100D8A82;
precomp_y[16] = 256'hB9C398F186806F5D27561506E4557433A2CF15009E498AE7ADEE9D63D01B2396;
precomp_y[17] = 256'h02972D2DE4F8D20681A78D93EC96FE23C26BFAE84FB14DB43B01E1E9056B8C49;
precomp_y[18] = 256'h80FC06BD8CC5B01098088A1950EED0DB01AA132967AB472235F5642483B25EAF;
precomp_y[19] = 256'h1C38303F1CC5C30F26E66BAD7FE72F70A65EED4CBE7024EB1AA01F56430BD57A;
precomp_y[20] = 256'h0D0E3FA9ECA8726909559E0D79269046BDC59EA10C70CE2B02D499EC224DC7F7;
precomp_y[21] = 256'hEECF41253136E5F99966F21881FD656EBC4345405C520DBC063465B521409933;
precomp_y[22] = 256'h758F3F41AFD6ED428B3081B0512FD62A54C3F3AFBB5B6764B653052A12949C9A;
precomp_y[23] = 256'h958EF42A7886B6400A08266E9BA1B37896C95330D97077CBBE8EB3C7671C60D6;
precomp_y[24] = 256'hE0DEDC9B3B2F8DAD4DA1F32DEC2531DF9EB5FBEB0598E4FD1A117DBA703A3C37;
precomp_y[25] = 256'h5ED430D78C296C3543114306DD8622D7C622E27C970A1DE31CB377B01AF7307E;
precomp_y[26] = 256'hCEDABD9B82203F7E13D206FCDF4E33D92A6C53C26E5CCE26D6579962C4E31DF6;
precomp_y[27] = 256'hCB474660EF35F5F2A41B643FA5E460575F4FA9B7962232A5C32F908318A04476;
precomp_y[28] = 256'h4119B88753C15BD6A693B03FCDDBB45D5AC6BE74AB5F0EF44B0BE9475A7E4B40;
precomp_y[29] = 256'h091B649609489D613D1D5E590F78E6D74ECFC061D57048BAD9E76F302C5B9C61;
precomp_y[30] = 256'h0673FB86E5BDA30FB3CD0ED304EA49A023EE33D0197A695D0C5D98093C536683;
precomp_y[31] = 256'h59C9E0BBA394E76F40C0AA58379A3CB6A5A2283993E90C4167002AF4920E37F5;
precomp_y[32] = 256'h3B952D32C67CF77E2E17446E204180AB21FB8090895138B4A4A797F86E80888B;
precomp_y[33] = 256'h55EB2DAFD84D6CCD5F862B785DC39D4AB157222720EF9DA217B8C45CF2BA2417;
precomp_y[34] = 256'hEFAE9C8DBC14130661E8CEC030C89AD0C13C66C0D17A2905CDC706AB7399A868;
precomp_y[35] = 256'hE38DA76DCD440621988D00BCF79AF25D5B29C094DB2A23146D003AFD41943E7A;
precomp_y[36] = 256'hF98A3FD831EB2B749A93B0E6F35CFB40C8CD5AA667A15581BC2FEDED498FD9C6;
precomp_y[37] = 256'h744B1152EACBE5E38DCC887980DA38B897584A65FA06CEDD2C924F97CBAC5996;
precomp_y[38] = 256'hC534AD44175FBC300F4EA6CE648309A042CE739A7919798CD85E216C4A307F6E;
precomp_y[39] = 256'hE13817B44EE14DE663BF4BC808341F326949E21A6A75C2570778419BDAF5733D;
precomp_y[40] = 256'h30E93E864E669D82224B967C3020B8FA8D1E4E350B6CBCC537A48B57841163A2;
precomp_y[41] = 256'hE491A42537F6E597D5D28A3224B1BC25DF9154EFBD2EF1D2CBBA2CAE5347D57E;
precomp_y[42] = 256'h100B610EC4FFB4760D5C1FC133EF6F6B12507A051F04AC5760AFA5B29DB83437;
precomp_y[43] = 256'hEF0AFBB2056205448E1652C48E8127FC6039E77C15C2378B7E7D15A0DE293311;
precomp_y[44] = 256'h8B378A22D827278D89C5E9BE8F9508AE3C2AD46290358630AFB34DB04EEDE0A4;
precomp_y[45] = 256'h68651CF9B6DA903E0914448C6CD9D4CA896878F5282BE4C8CC06E2A404078575;
precomp_y[46] = 256'hF5435A2BD2BADF7D485A4D8B8DB9FCCE3E1EF8E0201E4578C54673BC1DC5EA1D;
precomp_y[47] = 256'hD56EB30B69463E7234F5137B73B84177434800BACEBFC685FC37BBE9EFE4070D;
precomp_y[48] = 256'hEDD77F50BCB5A3CAB2E90737309667F2641462A54070F3D519212D39C197A629;
precomp_y[49] = 256'h0A855BABAD5CD60C88B430A69F53A1A7A38289154964799BE43D06D77D31DA06;
precomp_y[50] = 256'h66DB656F87D1F04FFFD1F04788C06830871EC5A64FEEE685BD80F0B1286D8374;
precomp_y[51] = 256'h09414685E97B1B5954BD46F730174136D57F1CEEB487443DC5321857BA73ABEE;
precomp_y[52] = 256'h4CB95957E83D40B0F73AF4544CCCF6B1F4B08D3C07B27FB8D8C2962A400766D1;
precomp_y[53] = 256'hFA77968128D9C92EE1010F337AD4717EFF15DB5ED3C049B3411E0315EAA4593B;
precomp_y[54] = 256'h5F3032F5892156E39CCD3D7915B9E1DA2E6DAC9E6F26E961118D14B8462E1661;
precomp_y[55] = 256'h8EC0BA238B96BEC0CBDDDCAE0AA442542EEE1FF50C986EA6B39847B3CC092FF6;
precomp_y[56] = 256'h8DC2412AAFE3BE5C4C5F37E0ECC5F9F6A446989AF04C4E25EBAAC479EC1C8C1E;
precomp_y[57] = 256'h5E4631150E62FB40D0E8C2A7CA5804A39D58186A50E497139626778E25B0674D;
precomp_y[58] = 256'hF65F5D3E292C2E0819A528391C994624D784869D7E6EA67FB18041024EDC07DC;
precomp_y[59] = 256'hF3E0319169EB9B85D5404795539A5E68FA1FBD583C064D2462B675F194A3DDB4;
precomp_y[60] = 256'h42242A969283A5F339BA7F075E36BA2AF925CE30D767ED6E55F4B031880D562C;
precomp_y[61] = 256'h204B5D6F84822C307E4B4A7140737AEC23FC63B65B35F86A10026DBD2D864E6B;
precomp_y[62] = 256'h04F14351D0087EFA49D245B328984989D5CAF9450F34BFC0ED16E96B58FA9913;
precomp_y[63] = 256'h073867F59C0659E81904F9A1C7543698E62562D6744C169CE7A36DE01A8D6154;
precomp_y[64] = 256'h39F23F366809085BEEBFC71181313775A99C9AED7D8BA38B161384C746012865;
precomp_y[65] = 256'hD2424B1B1ABE4EB8164227B085C9AA9456EA13493FD563E06FD51CF5694C78FC;
precomp_y[66] = 256'hEAD12168595FE1BE99252129B6E56B3391F7AB1410CD1E0EF3DCDCABD2FDA224;
precomp_y[67] = 256'h6FDCEF09F2F6D0A044E654AEF624136F503D459C3E89845858A47A9129CDD24E;
precomp_y[68] = 256'h060660257DD11B3AA9C8ED618D24EDFF2306D320F1D03010E33A7D2057F3B3B6;
precomp_y[69] = 256'h3D98A9CDD026DD43F39048F25A8847F4FCAFAD1895D7A633C6FED3C35E999511;
precomp_y[70] = 256'h0B4C4FE99C775A606E2D8862179139FFDA61DC861C019E55CD2876EB2A27D84B;
precomp_y[71] = 256'hAE434102EDDE0958EC4B19D917A6A28E6B72DA1834AFF0E650F049503A296CF2;
precomp_y[72] = 256'hCF2174118C8B6D7A4B48F6D534CE5C79422C086A63460502B827CE62A326683C;
precomp_y[73] = 256'h6FB8D5591B466F8FC63DB50F1C0F1C69013F996887B8244D2CDEC417AFEA8FA3;
precomp_y[74] = 256'h322AF4908C7312B0CFBFE369F7A7B3CDB7D4494BC2823700CFD652188A3EA98D;
precomp_y[75] = 256'h6749E67C029B85F52A034EAFD096836B2520818680E26AC8F3DFBCDB71749700;
precomp_y[76] = 256'h2AEABE7E4531510116217F07BF4D07300DE97E4874F81F533420A72EEB0BD6A4;
precomp_y[77] = 256'hB0EA558A113C30BEA60FC4775460C7901FF0B053D25CA2BDEEE98F1A4BE5D196;
precomp_y[78] = 256'h998C74A8CD45AC01289D5833A7BEB4744FF536B01B257BE4C5767BEA93EA57A4;
precomp_y[79] = 256'hB2284279995A34E2F9D4DE7396FC18B80F9B8B9FDD270F6661F79CA4C81BD257;
precomp_y[80] = 256'hBDD46039FEED17881D1E0862DB347F8CF395B74FC4BCDC4E940B74E3AC1F1B13;
precomp_y[81] = 256'h6F0A256BC5EFDF429A2FB6242F1A43A2D9B925BB4A4B3A26BB8E0F45EB596096;
precomp_y[82] = 256'hC359D6923BB398F7FD4473E16FE1C28475B740DD098075E6C0E8649113DC3A38;
precomp_y[83] = 256'h021AE7F4680E889BB130619E2C0F95A360CEB573C70603139862AFD617FA9B9F;
precomp_y[84] = 256'h60EA7F61A353524D1C987F6ECEC92F086D565AB687870CB12689FF1E31C74448;
precomp_y[85] = 256'h49B96715AB6878A79E78F07CE5680C5D6673051B4935BD897FEA824B77DC208A;
precomp_y[86] = 256'h5CA560753BE2A12FC6DE6CAF2CB489565DB936156B9514E1BB5E83037E0FA2D4;
precomp_y[87] = 256'h7571D74EE5E0FB92A7A8B33A07783341A5492144CC54BCC40A94473693606437;
precomp_y[88] = 256'hBE52D107BCFA09D8BCB9736A828CFA7FAC8DB17BF7A76A2C42AD961409018CF7;
precomp_y[89] = 256'h8FD64A14C06B589C26B947AE2BCF6BFA0149EF0BE14ED4D80F448A01C43B1C6D;
precomp_y[90] = 256'h39E5C9925B5A54B07433A4F18C61726F8BB131C012CA542EB24A8AC07200682A;
precomp_y[91] = 256'h62DFAF07A0F78FEB30E30D6295853CE189E127760AD6CF7FAE164E122A208D54;
precomp_y[92] = 256'h25A748AB367979D98733C38A1FA1C2E7DC6CC07DB2D60A9AE7A76AAA49BD0F77;
precomp_y[93] = 256'hECFB7056CF1DE042F9420BAB396793C0C390BDE74B4BBDFF16A83AE09A9A7517;
precomp_y[94] = 256'hCD450EC335438986DFEFA10C57FEA9BCC521A0959B2D80BBF74B190DCA712D10;
precomp_y[95] = 256'hF5C54754A8F71EE540B9B48728473E314F729AC5308B06938360990E2BFAD125;
precomp_y[96] = 256'h6CB9A8876D9CB8520609AF3ADD26CD20A0A7CD8A9411131CE85F44100099223E;
precomp_y[97] = 256'hFEF5A3C68059A6DEC5D624114BF1E91AAC2B9DA568D6ABEB2570D55646B8ADF1;
precomp_y[98] = 256'h1ACB250F255DD61C43D94CCC670D0F58F49AE3FA15B96623E5430DA0AD6C62B2;
precomp_y[99] = 256'h5F310D4B3C99B9EBB19F77D41C1DEE018CF0D34FD4191614003E945A1216E423;
precomp_y[100] = 256'h438136D603E858A3A5C440C38ECCBADDC1D2942114E2EDDD4740D098CED1F0D8;
precomp_y[101] = 256'hCDB559EEDC2D79F926BAF44FB84EA4D44BCF50FEE51D7CEB30E2E7F463036758;
precomp_y[102] = 256'h0C3B997D050EE5D423EBAF66A6DB9F57B3180C902875679DE924B69D84A7B375;
precomp_y[103] = 256'h6D89AD7BA4876B0B22C2CA280C682862F342C8591F1DAF5170E07BFD9CCAFA7D;
precomp_y[104] = 256'hCA5EF7D4B231C94C3B15389A5F6311E9DAFF7BB67B103E9880EF4BFF637ACAEC;
precomp_y[105] = 256'h09731141D81FC8F8084D37C6E7542006B3EE1B40D60DFE5362A5B132FD17DDC0;
precomp_y[106] = 256'hEE1849F513DF71E32EFC3896EE28260C73BB80547AE2275BA497237794C8753C;
precomp_y[107] = 256'hD3AA2ED71C9DD2247A62DF062736EB0BADDEA9E36122D2BE8641ABCB005CC4A4;
precomp_y[108] = 256'hC4E1020916980A4DA5D01AC5E6AD330734EF0D7906631C4F2390426B2EDD791F;
precomp_y[109] = 256'h67163E903236289F776F22C25FB8A3AFC1732F2B84B4E95DBDA47AE5A0852649;
precomp_y[110] = 256'h0CD1BC7CB6CC407BB2F0CA647C718A730CF71872E7D0D2A53FA20EFCDFE61826;
precomp_y[111] = 256'h299D21F9413F33B3EDF43B257004580B70DB57DA0B182259E09EECC69E0D38A5;
precomp_y[112] = 256'hF9429E738B8E53B968E99016C059707782E14F4535359D582FC416910B3EEA87;
precomp_y[113] = 256'h462F9BCE619898638499350113BBC9B10A878D35DA70740DC695A559EB88DB7B;
precomp_y[114] = 256'h62188BC49D61E5428573D48A74E1C655B1C61090905682A0D5558ED72DCCB9BC;
precomp_y[115] = 256'h7C10DFB164C3425F5C71A3F9D7992038F1065224F72BB9D1D902A6D13037B47C;
precomp_y[116] = 256'hAB8C1E086D04E813744A655B2DF8D5F83B3CDC6FAA3088C1D3AEA1454E3A1D5F;
precomp_y[117] = 256'h4CB04437F391ED73111A13CC1D4DD0DB1693465C2240480D8955E8592F27447A;
precomp_y[118] = 256'hBD1AEB21AD22EBB22A10F0303417C6D964F8CDD7DF0ACA614B10DC14D125AC46;
precomp_y[119] = 256'hBFEFACDB0E5D0FD7DF3A311A94DE062B26B80C61FBC97508B79992671EF7CA7F;
precomp_y[120] = 256'h603C12DAF3D9862EF2B25FE1DE289AED24ED291E0EC6708703A5BD567F32ED03;
precomp_y[121] = 256'hCC6157EF18C9C63CD6193D83631BBEA0093E0968942E8C33D5737FD790E0DB08;
precomp_y[122] = 256'h553E04F6B018B4FA6C8F39E7F311D3176290D0E0F19CA73F17714D9977A22FF8;
precomp_y[123] = 256'h0712FCDD1B9053F09003A3481FA7762E9FFD7C8EF35A38509E2FBF2629008373;
precomp_y[124] = 256'hED8CC9D04B29EB877D270B4878DC43C19AEFD31F4EEE09EE7B47834C1FA4B1C3;
precomp_y[125] = 256'h9852390A99507679FD0B86FD2B39A868D7EFC22151346E1A3CA4726586A6BED8;
precomp_y[126] = 256'h9E994980D9917E22B76B061927FA04143D096CCC54963E6A5EBFA5F3F8E286C1;
precomp_y[127] = 256'h4036EDC931A60AE889353F77FD53DE4A2708B26B6F5DA72AD3394119DAF408F9;
