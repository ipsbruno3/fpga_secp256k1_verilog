precomp_y[0] = 256'h483ADA7726A3C4655DA4FBFC0E1108A8FD17B448A68554199C47D08FFB10D4B8;
precomp_y[1] = 256'h388F7B0F632DE8140FE337E62A37F3566500A99934C2231B6CB9FD7584B8E672;
precomp_y[2] = 256'hD8AC222636E5E3D6D4DBA9DDA6C9C426F788271BAB0D6840DCA87D3AA6AC62D6;
precomp_y[3] = 256'h6AEBCA40BA255960A3178D6D861A54DBA813D0B813FDE7B5A5082628087264DA;
precomp_y[4] = 256'hCC338921B0A7D9FD64380971763B61E9ADD888A4375F8E0F05CC262AC64F9C37;
precomp_y[5] = 256'hD984A032EB6B5E190243DD56D7B7B365372DB1E2DFF9D6A8301D74C9C953C61B;
precomp_y[6] = 256'h0AB0902E8D880A89758212EB65CDAF473A1A06DA521FA91F29B5CB52DB03ED81;
precomp_y[7] = 256'h581E2872A86C72A683842EC228CC6DEFEA40AF2BD896D3A5C504DC9FF6A26B58;
precomp_x[0] = 256'h79BE667EF9DCBBAC55A06295CE870B07029BFCDB2DCE28D959F2815B16F81798;
precomp_x[1] = 256'hF9308A019258C31049344F85F89D5229B531C845836F99B08601F113BCE036F9;
precomp_x[2] = 256'h2F8BDE4D1A07209355B4A7250A5C5128E88B84BDDC619AB7CBA8D569B240EFE4;
precomp_x[3] = 256'h5CBDF0646E5DB4EAA398F365F2EA7A0E3D419B7E0330E39CE92BDDEDCAC4F9BC;
precomp_x[4] = 256'hACD484E2F0C7F65309AD178A9F559ABDE09796974C57E714C35F110DFC27CCBE;
precomp_x[5] = 256'h774AE7F858A9411E5EF4246B70C65AAC5649980BE5C17891BBEC17895DA008CB;
precomp_x[6] = 256'hF28773C2D975288BC7D1D205C3748651B075FBC6610E58CDDEEDDF8F19405AA8;
precomp_x[7] = 256'hD7924D4F7D43EA965A465AE3095FF41131E5946F3C85F79E44ADBCF8E27E080E;
